magic
tech sky130A
magscale 1 2
timestamp 1726787590
<< nwell >>
rect -920 920 -400 960
rect -920 420 -880 920
rect -760 760 -560 860
rect -543 760 -509 776
rect -820 740 -811 760
rect -777 740 -500 760
rect -820 600 -500 740
rect -820 580 -811 600
rect -777 580 -500 600
rect -760 480 -560 580
rect -543 574 -509 580
rect -440 420 -400 920
rect -920 380 -400 420
<< nbase >>
rect -960 960 -360 1000
rect -960 380 -920 960
rect -880 860 -440 920
rect -880 760 -760 860
rect -560 776 -440 860
rect -560 760 -543 776
rect -509 760 -440 776
rect -880 580 -820 760
rect -811 740 -777 760
rect -811 580 -777 600
rect -500 580 -440 760
rect -880 480 -760 580
rect -560 574 -543 580
rect -509 574 -440 580
rect -560 480 -440 574
rect -880 420 -440 480
rect -400 380 -360 960
rect -960 340 -360 380
<< pmos >>
rect -760 580 -560 760
<< pdiff >>
rect -820 740 -760 760
rect -820 600 -811 740
rect -777 600 -760 740
rect -820 580 -760 600
rect -560 740 -500 760
rect -560 600 -543 740
rect -509 600 -500 740
rect -560 580 -500 600
<< pdiffc >>
rect -811 600 -777 740
rect -543 600 -509 740
<< nsubdiff >>
rect -920 920 -820 960
rect -500 920 -400 960
rect -920 840 -880 920
rect -440 840 -400 920
rect -920 420 -880 480
rect -440 420 -400 480
rect -920 380 -820 420
rect -500 380 -400 420
<< nsubdiffcont >>
rect -820 920 -500 960
rect -920 480 -880 840
rect -440 480 -400 840
rect -820 380 -500 420
<< poly >>
rect -760 844 -560 860
rect -760 810 -740 844
rect -580 810 -560 844
rect -760 760 -560 810
rect -760 529 -560 580
rect -760 495 -740 529
rect -580 495 -560 529
rect -760 480 -560 495
<< polycont >>
rect -740 810 -580 844
rect -740 495 -580 529
<< locali >>
rect -920 920 -820 960
rect -500 920 -400 960
rect -920 840 -880 920
rect -760 810 -740 844
rect -580 810 -560 844
rect -440 840 -400 920
rect -811 740 -777 775
rect -811 567 -777 600
rect -543 740 -509 776
rect -543 568 -509 600
rect -760 495 -740 529
rect -580 495 -560 529
rect -920 420 -880 480
rect -440 420 -400 480
rect -920 380 -820 420
rect -500 380 -400 420
<< viali >>
rect -740 810 -580 844
rect -811 600 -777 740
rect -543 600 -509 740
rect -740 495 -580 529
<< metal1 >>
rect -752 844 -568 856
rect -752 840 -740 844
rect -760 810 -740 840
rect -580 840 -568 844
rect -580 810 -560 840
rect -752 800 -568 810
rect -818 740 -770 760
rect -818 600 -811 740
rect -777 600 -770 740
rect -818 580 -770 600
rect -550 740 -502 760
rect -550 600 -543 740
rect -509 600 -502 740
rect -550 580 -502 600
rect -753 529 -567 541
rect -753 495 -740 529
rect -580 495 -567 529
rect -753 483 -567 495
<< labels >>
flabel nsubdiffcont -660 940 -660 940 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel viali -660 820 -660 820 0 FreeSans 400 0 0 0 G
port 1 nsew
flabel viali -800 680 -800 680 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel viali -520 680 -520 680 0 FreeSans 400 0 0 0 D
port 0 nsew
<< end >>
