magic
tech sky130A
timestamp 1730605901
<< nwell >>
rect -344 -1031 344 1031
<< pmos >>
rect -297 -1000 -247 1000
rect -161 -1000 -111 1000
rect -25 -1000 25 1000
rect 111 -1000 161 1000
rect 247 -1000 297 1000
<< pdiff >>
rect -326 994 -297 1000
rect -326 -994 -320 994
rect -303 -994 -297 994
rect -326 -1000 -297 -994
rect -247 994 -218 1000
rect -247 -994 -241 994
rect -224 -994 -218 994
rect -247 -1000 -218 -994
rect -190 994 -161 1000
rect -190 -994 -184 994
rect -167 -994 -161 994
rect -190 -1000 -161 -994
rect -111 994 -82 1000
rect -111 -994 -105 994
rect -88 -994 -82 994
rect -111 -1000 -82 -994
rect -54 994 -25 1000
rect -54 -994 -48 994
rect -31 -994 -25 994
rect -54 -1000 -25 -994
rect 25 994 54 1000
rect 25 -994 31 994
rect 48 -994 54 994
rect 25 -1000 54 -994
rect 82 994 111 1000
rect 82 -994 88 994
rect 105 -994 111 994
rect 82 -1000 111 -994
rect 161 994 190 1000
rect 161 -994 167 994
rect 184 -994 190 994
rect 161 -1000 190 -994
rect 218 994 247 1000
rect 218 -994 224 994
rect 241 -994 247 994
rect 218 -1000 247 -994
rect 297 994 326 1000
rect 297 -994 303 994
rect 320 -994 326 994
rect 297 -1000 326 -994
<< pdiffc >>
rect -320 -994 -303 994
rect -241 -994 -224 994
rect -184 -994 -167 994
rect -105 -994 -88 994
rect -48 -994 -31 994
rect 31 -994 48 994
rect 88 -994 105 994
rect 167 -994 184 994
rect 224 -994 241 994
rect 303 -994 320 994
<< poly >>
rect -297 1000 -247 1013
rect -161 1000 -111 1013
rect -25 1000 25 1013
rect 111 1000 161 1013
rect 247 1000 297 1013
rect -297 -1013 -247 -1000
rect -161 -1013 -111 -1000
rect -25 -1013 25 -1000
rect 111 -1013 161 -1000
rect 247 -1013 297 -1000
<< locali >>
rect -320 994 -303 1002
rect -320 -1002 -303 -994
rect -241 994 -224 1002
rect -241 -1002 -224 -994
rect -184 994 -167 1002
rect -184 -1002 -167 -994
rect -105 994 -88 1002
rect -105 -1002 -88 -994
rect -48 994 -31 1002
rect -48 -1002 -31 -994
rect 31 994 48 1002
rect 31 -1002 48 -994
rect 88 994 105 1002
rect 88 -1002 105 -994
rect 167 994 184 1002
rect 167 -1002 184 -994
rect 224 994 241 1002
rect 224 -1002 241 -994
rect 303 994 320 1002
rect 303 -1002 320 -994
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l .5 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_01v8_S2VXMU parameters
<< end >>
