magic
tech sky130A
magscale 1 2
timestamp 1733331218
<< nwell >>
rect 9000 -11600 29200 1400
<< pwell >>
rect 3800 1400 32200 3600
rect 3800 -11600 9000 1400
rect 29200 -1034 32200 1400
rect 29200 -2840 30124 -1034
rect 31970 -2840 32200 -1034
rect 29200 -11600 32200 -2840
rect 3800 -12000 32200 -11600
<< psubdiff >>
rect 3800 3550 32200 3600
rect 3800 3450 4200 3550
rect 31600 3450 32200 3550
rect 3800 3400 32200 3450
rect 3800 3250 4000 3400
rect 3800 -11450 3850 3250
rect 3950 -11450 4000 3250
rect 32000 3250 32200 3400
rect 3800 -11800 4000 -11450
rect 32000 -11700 32050 3250
rect 32150 -11700 32200 3250
rect 32000 -11800 32200 -11700
rect 3800 -11850 32200 -11800
rect 3800 -11950 4200 -11850
rect 31850 -11950 32200 -11850
rect 3800 -12000 32200 -11950
<< nsubdiff >>
rect 9200 1150 29100 1200
rect 9200 1050 10350 1150
rect 28500 1050 29100 1150
rect 9200 1000 29100 1050
rect 9200 -10950 9250 1000
rect 9350 -10950 9400 1000
rect 9200 -11300 9400 -10950
rect 28900 250 29100 1000
rect 28900 -10850 28950 250
rect 29050 -10850 29100 250
rect 28900 -11300 29100 -10850
rect 9200 -11350 29100 -11300
rect 9200 -11450 9750 -11350
rect 28400 -11450 29100 -11350
rect 9200 -11500 29100 -11450
<< psubdiffcont >>
rect 4200 3450 31600 3550
rect 3850 -11450 3950 3250
rect 32050 -11700 32150 3250
rect 4200 -11950 31850 -11850
<< nsubdiffcont >>
rect 10350 1050 28500 1150
rect 9250 -10950 9350 1000
rect 28950 -10850 29050 250
rect 9750 -11450 28400 -11350
<< locali >>
rect 3800 3550 32200 3600
rect 3800 3450 4200 3550
rect 31600 3450 32200 3550
rect 3800 3400 32200 3450
rect 3800 3250 5504 3400
rect 3800 -11450 3850 3250
rect 3950 1500 5504 3250
rect 32000 3250 32200 3400
rect 3950 1350 5600 1500
rect 3950 -520 4000 1350
rect 9200 1150 29100 1200
rect 5596 1072 5600 1100
rect 5020 960 5600 1072
rect 9200 1050 10350 1150
rect 28500 1050 29100 1150
rect 9200 1000 29100 1050
rect 4320 180 4600 220
rect 4320 -100 4340 180
rect 4380 160 4600 180
rect 4380 -100 4560 160
rect 4320 -160 4560 -100
rect 4320 -180 4600 -160
rect 8160 -260 8520 160
rect 3950 -940 4400 -520
rect 3950 -3150 4000 -940
rect 4800 -1260 5000 -1200
rect 7800 -1240 8000 -1200
rect 4800 -1600 4920 -1260
rect 7900 -1300 8000 -1240
rect 7900 -1360 7920 -1300
rect 7980 -1360 8000 -1300
rect 7900 -1600 8000 -1360
rect 8460 -2720 8520 -760
rect 8460 -2800 8480 -2720
rect 5260 -2876 5820 -2800
rect 8460 -2820 8520 -2800
rect 3950 -3168 5258 -3150
rect 5834 -3168 5850 -3150
rect 3950 -3200 5850 -3168
rect 3950 -3240 8480 -3200
rect 8520 -3240 8900 -3200
rect 3950 -11450 8900 -3240
rect 3800 -11800 8900 -11450
rect 9200 -10950 9250 1000
rect 9350 -10950 9400 1000
rect 28900 250 29100 1000
rect 21000 -240 21040 -200
rect 21000 -260 21200 -240
rect 12400 -1000 13400 -800
rect 10000 -1200 13400 -1000
rect 10000 -1460 10200 -1200
rect 10000 -1540 10060 -1460
rect 10140 -1540 10200 -1460
rect 10000 -1800 10200 -1540
rect 9200 -11300 9400 -10950
rect 28900 -10850 28950 250
rect 29050 -10850 29100 250
rect 32000 -600 32050 3250
rect 29550 -950 32050 -600
rect 32000 -2700 32050 -950
rect 31998 -2914 32050 -2700
rect 28900 -11300 29100 -10850
rect 9200 -11350 29100 -11300
rect 9200 -11450 9750 -11350
rect 28400 -11450 29100 -11350
rect 9200 -11500 29100 -11450
rect 29300 -4650 32050 -2914
rect 29300 -4750 29600 -4650
rect 29750 -4750 32050 -4650
rect 29300 -11700 32050 -4750
rect 32150 -11700 32200 3250
rect 29300 -11800 32200 -11700
rect 3800 -11850 32200 -11800
rect 3800 -11950 4200 -11850
rect 31850 -11950 32200 -11850
rect 3800 -12000 32200 -11950
<< viali >>
rect 9560 1840 9760 1960
rect 5644 1134 5678 1302
rect 5018 1072 5594 1106
rect 10350 1050 28500 1150
rect 5660 860 5860 940
rect 4330 540 4380 680
rect 8480 530 8520 630
rect 4340 -100 4380 180
rect 4560 -160 4620 160
rect 5900 -1160 6100 -1040
rect 7920 -1360 7980 -1300
rect 5280 -1540 5360 -1480
rect 7380 -1540 7560 -1460
rect 8480 -2800 8520 -2720
rect 5258 -2910 5834 -2876
rect 5884 -3106 5918 -2938
rect 5258 -3168 5834 -3134
rect 8480 -3240 8520 -3200
rect 10440 460 13600 500
rect 20640 440 21560 560
rect 25180 540 26300 660
rect 17420 -240 17560 -200
rect 21040 -240 21200 -200
rect 10860 -740 11360 -660
rect 25960 -1460 26180 -1360
rect 28040 -1460 28230 -1350
rect 10060 -1540 10140 -1460
rect 26660 -4820 26700 -4700
rect 29344 -556 29512 -522
rect 29282 -982 29316 -606
rect 30342 -1919 30376 -1885
rect 29600 -4750 29750 -4650
<< metal1 >>
rect 3800 3400 32200 3600
rect 3800 1496 5504 3400
rect 5640 3000 29500 3200
rect 3800 -11800 4000 1496
rect 5640 1302 5680 3000
rect 5640 1140 5644 1302
rect 5678 1140 5680 1302
rect 5540 940 5960 960
rect 5540 860 5660 940
rect 5860 860 5960 940
rect 5540 840 5960 860
rect 4320 680 4400 700
rect 4320 540 4330 680
rect 4390 540 4400 680
rect 4320 520 4400 540
rect 8460 630 8540 650
rect 8520 530 8540 630
rect 8460 510 8540 530
rect 4220 180 4640 200
rect 4220 -100 4340 180
rect 4380 160 4640 180
rect 4380 -100 4560 160
rect 4220 -160 4560 -100
rect 4620 -160 4640 160
rect 4220 -180 4640 -160
rect 5860 -1040 6140 -1000
rect 5860 -1160 5900 -1040
rect 6100 -1160 6140 -1040
rect 5860 -1200 6140 -1160
rect 7900 -1300 8000 -1280
rect 7900 -1360 7920 -1300
rect 7980 -1360 8000 -1300
rect 7900 -1380 8000 -1360
rect 7360 -1460 7580 -1440
rect 5240 -1480 5400 -1460
rect 5240 -1540 5280 -1480
rect 5360 -1540 5400 -1480
rect 5240 -1560 5400 -1540
rect 7360 -1540 7380 -1460
rect 7560 -1540 7580 -1460
rect 7360 -1580 7580 -1540
rect 8460 -2700 8520 -760
rect 8440 -2720 8540 -2700
rect 8440 -2800 8460 -2720
rect 8520 -2800 8540 -2720
rect 8440 -2840 8540 -2800
rect 5880 -3080 5884 -2940
rect 8600 -2940 8800 3000
rect 9400 1960 28560 2800
rect 9400 1840 9560 1960
rect 9760 1840 28560 1960
rect 9400 1150 28560 1840
rect 9400 1050 10350 1150
rect 28500 1050 28560 1150
rect 9400 660 28560 1050
rect 9400 600 25180 660
rect 10420 500 13620 600
rect 10420 460 10440 500
rect 13600 460 13620 500
rect 10420 440 13620 460
rect 20400 560 21600 600
rect 20400 440 20640 560
rect 21560 440 21600 560
rect 24480 540 25180 600
rect 26300 540 28560 660
rect 24480 500 28560 540
rect 20400 400 21600 440
rect 17400 -200 17580 -180
rect 17400 -260 17420 -200
rect 17560 -260 17580 -200
rect 21000 -200 21220 -180
rect 21000 -220 21040 -200
rect 17400 -280 17580 -260
rect 21020 -280 21040 -220
rect 21200 -280 21220 -200
rect 21020 -300 21220 -280
rect 29400 -522 29500 3000
rect 29400 -580 29500 -556
rect 10820 -660 11380 -640
rect 10820 -740 10860 -660
rect 11360 -740 11380 -660
rect 10820 -760 11380 -740
rect 29250 -720 29282 -710
rect 29250 -850 29282 -840
rect 29316 -850 29320 -710
rect 30260 -1158 30866 -1156
rect 30260 -1190 31832 -1158
rect 25900 -1360 26240 -1340
rect 10040 -1460 10160 -1440
rect 10040 -1540 10060 -1460
rect 10140 -1540 10160 -1460
rect 25900 -1460 25960 -1360
rect 26180 -1460 26240 -1360
rect 25900 -1480 26240 -1460
rect 28010 -1350 28280 -1310
rect 28010 -1460 28040 -1350
rect 28230 -1460 28280 -1350
rect 28010 -1500 28280 -1460
rect 10040 -1560 10160 -1540
rect 30260 -1714 31836 -1190
rect 30260 -1872 30866 -1714
rect 30260 -1926 30334 -1872
rect 30386 -1926 30866 -1872
rect 30260 -2160 30866 -1926
rect 30977 -2023 31147 -1853
rect 31246 -2160 31836 -1714
rect 30258 -2724 31836 -2160
rect 30258 -2726 31816 -2724
rect 30260 -2736 30866 -2726
rect 5918 -3080 8800 -2940
rect 8460 -3180 8560 -3160
rect 8460 -3240 8480 -3180
rect 8540 -3240 8560 -3180
rect 8460 -3260 8560 -3240
rect 29550 -4650 29800 -4600
rect 26640 -4700 26720 -4680
rect 26640 -4820 26660 -4700
rect 29550 -4750 29600 -4650
rect 29750 -4750 29800 -4650
rect 29550 -4800 29800 -4750
rect 26640 -4840 26720 -4820
rect 32000 -11800 32200 3400
rect 3800 -12000 32200 -11800
<< via1 >>
rect 4330 540 4380 680
rect 4380 540 4390 680
rect 8460 530 8480 630
rect 8480 530 8520 630
rect 5900 -1160 6100 -1040
rect 7920 -1360 7980 -1300
rect 5280 -1540 5360 -1480
rect 7380 -1540 7560 -1460
rect 8460 -2800 8480 -2720
rect 8480 -2800 8520 -2720
rect 9560 1840 9760 1960
rect 17420 -240 17560 -200
rect 17420 -260 17560 -240
rect 21040 -240 21200 -200
rect 21040 -280 21200 -240
rect 10860 -740 11360 -660
rect 29250 -840 29282 -720
rect 29282 -840 29310 -720
rect 10060 -1540 10140 -1460
rect 25960 -1460 26180 -1360
rect 28040 -1460 28230 -1350
rect 30334 -1885 30386 -1872
rect 30334 -1919 30342 -1885
rect 30342 -1919 30376 -1885
rect 30376 -1919 30386 -1885
rect 30334 -1926 30386 -1919
rect 8480 -3200 8540 -3180
rect 8480 -3240 8520 -3200
rect 8520 -3240 8540 -3200
rect 26660 -4820 26700 -4700
rect 26700 -4820 26720 -4700
rect 29600 -4750 29750 -4650
<< metal2 >>
rect 8400 1960 9800 2000
rect 8400 1840 9560 1960
rect 9760 1840 9800 1960
rect 8400 1800 9800 1840
rect 4320 680 4400 700
rect 4320 540 4330 680
rect 4390 650 4400 680
rect 8400 650 8600 1800
rect 4390 630 8600 650
rect 4390 540 8460 630
rect 4320 530 8460 540
rect 8520 600 8600 630
rect 8520 530 8540 600
rect 4320 520 8540 530
rect 8460 510 8540 520
rect 17400 -200 17580 -180
rect 21000 -200 21220 -180
rect 17400 -260 17420 -200
rect 17560 -260 17600 -200
rect 10820 -660 11380 -640
rect 10820 -700 10860 -660
rect 5200 -740 10860 -700
rect 11360 -700 11380 -660
rect 11360 -740 11400 -700
rect 5200 -800 11400 -740
rect 5200 -1480 5400 -800
rect 17400 -1000 17600 -260
rect 5800 -1040 17600 -1000
rect 5800 -1160 5900 -1040
rect 6100 -1160 17600 -1040
rect 5800 -1200 17600 -1160
rect 21000 -280 21040 -200
rect 21200 -280 21220 -200
rect 21000 -1280 21220 -280
rect 7900 -1300 21220 -1280
rect 7900 -1360 7920 -1300
rect 7980 -1360 21220 -1300
rect 29200 -710 29300 -600
rect 29200 -720 29320 -710
rect 29200 -840 29250 -720
rect 29310 -840 29320 -720
rect 29200 -850 29320 -840
rect 7900 -1380 21220 -1360
rect 25900 -1360 26240 -1340
rect 5200 -1540 5280 -1480
rect 5360 -1540 5400 -1480
rect 5200 -1600 5400 -1540
rect 7360 -1460 10160 -1440
rect 7360 -1540 7380 -1460
rect 7560 -1540 10060 -1460
rect 10140 -1540 10160 -1460
rect 25900 -1460 25960 -1360
rect 26180 -1460 26240 -1360
rect 25900 -1480 26240 -1460
rect 28010 -1350 28280 -1310
rect 28010 -1460 28040 -1350
rect 28230 -1400 28280 -1350
rect 29200 -1400 29300 -850
rect 28230 -1460 29300 -1400
rect 7360 -1560 10160 -1540
rect 7360 -1580 7580 -1560
rect 26000 -1800 26200 -1480
rect 28010 -1500 29300 -1460
rect 26000 -1872 30400 -1800
rect 26000 -1926 30334 -1872
rect 30386 -1926 30400 -1872
rect 26000 -2000 30400 -1926
rect 8440 -2720 8540 -2700
rect 8440 -2800 8460 -2720
rect 8520 -2800 8540 -2720
rect 8440 -2840 8540 -2800
rect 8460 -3160 8540 -2840
rect 8460 -3180 8560 -3160
rect 8460 -3240 8480 -3180
rect 8540 -3240 8560 -3180
rect 8460 -3260 8560 -3240
rect 26700 -4650 29800 -4600
rect 26700 -4680 29600 -4650
rect 26640 -4700 29600 -4680
rect 26640 -4820 26660 -4700
rect 26720 -4750 29600 -4700
rect 29750 -4750 29800 -4650
rect 26720 -4800 29800 -4750
rect 26640 -4840 26720 -4820
use diff80  diff80_0
timestamp 1732736100
transform 1 0 20560 0 1 -300
box -3560 0 3800 840
use n1x15_diff_pair  n1x15_diff_pair_0
timestamp 1732735151
transform 1 0 5960 0 1 -1680
box -1360 -1320 2300 480
use n1x30_diff_pair  n1x30_diff_pair_0
timestamp 1732735011
transform 1 0 5760 0 -1 -1040
box -1360 -2240 2700 360
use p1_80x80  p1_80x80_0
timestamp 1732734633
transform 1 0 20820 0 -1 -11380
box -10800 -9960 6000 -120
use p1x15_diif_pair  p1x15_diif_pair_0
timestamp 1732735194
transform 1 0 11280 0 1 240
box -1080 -1240 2520 560
use p1x30_diff_pair  p1x30_diff_pair_0
timestamp 1732735234
transform 1 0 25860 0 1 380
box -1120 -2080 2880 520
use sky130_fd_pr__nfet_01v8_Q7B869  sky130_fd_pr__nfet_01v8_Q7B869_0
timestamp 1732757215
transform 1 0 29428 0 -1 -763
box -158 -257 158 257
use sky130_fd_pr__nfet_01v8_QX2DR5  sky130_fd_pr__nfet_01v8_QX2DR5_0
timestamp 1733160839
transform 0 1 5337 -1 0 1218
box -158 -357 158 357
use sky130_fd_pr__nfet_01v8_QX2DR5  sky130_fd_pr__nfet_01v8_QX2DR5_1
timestamp 1733160839
transform 0 1 5577 -1 0 -3022
box -158 -357 158 357
use sky130_fd_pr__res_xhigh_po_0p35_AS6SD6  sky130_fd_pr__res_xhigh_po_0p35_AS6SD6_0
timestamp 1732738914
transform 1 0 1300 0 1 -13500
box 0 0 1 1
use sky130_fd_pr__res_xhigh_po_0p35_AS6UD6  sky130_fd_pr__res_xhigh_po_0p35_AS6UD6_0
timestamp 1732738914
transform 1 0 1300 0 1 -13500
box 0 0 1 1
use sky130_fd_pr__res_xhigh_po_0p35_FPZZTN  sky130_fd_pr__res_xhigh_po_0p35_FPZZTN_0
timestamp 1732738914
transform 1 0 2750 0 1 1600
box 0 0 1 1
use sky130_fd_pr__res_xhigh_po_0p35_V22KJH  sky130_fd_pr__res_xhigh_po_0p35_V22KJH_0
timestamp 1732758882
transform 1 0 4355 0 1 -349
box -35 -591 35 591
use sky130_fd_pr__res_xhigh_po_0p35_V22KJH  sky130_fd_pr__res_xhigh_po_0p35_V22KJH_1
timestamp 1732758882
transform 1 0 8495 0 1 -429
box -35 -591 35 591
use sky130_fd_pr__res_xhigh_po_0p35_Y6F53N  sky130_fd_pr__res_xhigh_po_0p35_Y6F53N_0
timestamp 1732758882
transform 1 0 4355 0 1 306
box -35 -486 35 486
use sky130_fd_pr__res_xhigh_po_0p35_Y6F53N  sky130_fd_pr__res_xhigh_po_0p35_Y6F53N_1
timestamp 1732758882
transform 1 0 8495 0 1 226
box -35 -486 35 486
use sky130_fd_pr__rf_npn_05v5_W1p00L1p00  sky130_fd_pr__rf_npn_05v5_W1p00L1p00_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704896540
transform 1 0 30200 0 1 -2800
box 0 0 1724 1724
<< labels >>
flabel locali 8500 -20 8500 -20 0 FreeSans 1600 0 0 0 Vinn
flabel via1 6000 -1100 6000 -1100 0 FreeSans 1600 0 0 0 Vp
flabel via1 10100 -1500 10100 -1500 0 FreeSans 1600 0 0 0 Vg
flabel nwell 27740 -1390 27740 -1390 0 FreeSans 1600 0 0 0 Vd
flabel metal1 17160 2140 17160 2140 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 4270 60 4270 60 0 FreeSans 1600 0 0 0 Vinp
port 2 nsew
flabel pwell 6420 -2700 6420 -2700 0 FreeSans 1600 0 0 0 Vdiff2
flabel pwell 5760 900 5760 900 0 FreeSans 1600 0 0 0 Vdiff
flabel metal1 8706 3086 8706 3086 0 FreeSans 1600 0 0 0 Vref
port 4 nsew
flabel pwell 4616 2952 4616 2952 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel via1 30356 -1904 30356 -1904 0 FreeSans 1600 0 0 0 Vdo
flabel metal1 31062 -1936 31062 -1936 0 FreeSans 1600 0 0 0 Vout
port 5 nsew
<< properties >>
string demod parameters
<< end >>
