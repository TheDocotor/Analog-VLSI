magic
tech sky130A
magscale 1 2
timestamp 1729279979
use sky130_fd_pr__res_xhigh_po_0p69_2LTKQM  sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_0
timestamp 1729279979
transform 1 0 727 0 1 393
box -69 -761 69 761
use sky130_fd_pr__res_xhigh_po_0p69_2LTKQM  sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1
timestamp 1729279979
transform 1 0 729 0 1 -699
box -69 -761 69 761
<< end >>
