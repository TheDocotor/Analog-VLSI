magic
tech sky130A
timestamp 1726503206
<< error_p >>
rect -1022 1055 -577 1057
<< pwell >>
rect -1153 -49 -454 1146
<< nmos >>
rect -1040 52 -565 1038
<< ndiff >>
rect -1067 52 -1040 1038
rect -565 52 -537 1038
<< poly >>
rect -1040 1072 -565 1077
rect -1040 1055 -1022 1072
rect -577 1055 -565 1072
rect -1040 1038 -565 1055
rect -1040 33 -565 52
rect -1040 16 -1022 33
rect -577 16 -565 33
rect -1040 5 -565 16
<< polycont >>
rect -1022 1055 -577 1072
rect -1022 16 -577 33
<< locali >>
rect -1131 1122 -473 1124
rect -1133 1101 -473 1122
rect -1133 -13 -1111 1101
rect -1040 1055 -1022 1072
rect -577 1055 -565 1072
rect -1060 52 -1043 1038
rect -560 52 -540 1038
rect -1040 16 -1022 33
rect -577 16 -565 33
rect -490 -13 -473 1101
rect -1133 -30 -473 -13
<< viali >>
rect -1022 1055 -577 1072
rect -1022 16 -577 33
<< metal1 >>
rect -1036 1072 -570 1075
rect -1036 1055 -1022 1072
rect -577 1055 -570 1072
rect -1036 1050 -570 1055
rect -1032 33 -570 38
rect -1032 16 -1022 33
rect -577 16 -570 33
rect -1032 13 -570 16
use sky130_fd_pr__nfet_01v8_TSEK3K  sky130_fd_pr__nfet_01v8_TSEK3K_0
timestamp 1726503206
transform 1 0 811 0 1 902
box -348 -605 348 605
<< end >>
