magic
tech sky130A
magscale 1 2
timestamp 1728490836
<< pwell >>
rect -1400 200 0 2600
<< nmos >>
rect -1220 400 -1000 2400
rect -940 400 -720 2400
rect -660 400 -440 2400
rect -380 400 -160 2400
<< ndiff >>
rect -1280 2380 -1220 2400
rect -1280 420 -1265 2380
rect -1231 420 -1220 2380
rect -1280 400 -1220 420
rect -1000 2380 -940 2400
rect -1000 420 -985 2380
rect -951 420 -940 2380
rect -1000 400 -940 420
rect -720 2380 -660 2400
rect -720 420 -705 2380
rect -671 420 -660 2380
rect -720 400 -660 420
rect -440 2380 -380 2400
rect -440 420 -425 2380
rect -391 420 -380 2380
rect -440 400 -380 420
rect -160 2380 -100 2400
rect -160 420 -145 2380
rect -111 420 -100 2380
rect -160 400 -100 420
<< ndiffc >>
rect -1265 420 -1231 2380
rect -985 420 -951 2380
rect -705 420 -671 2380
rect -425 420 -391 2380
rect -145 420 -111 2380
<< poly >>
rect -1220 2480 -1000 2500
rect -1220 2440 -1200 2480
rect -1020 2440 -1000 2480
rect -1220 2400 -1000 2440
rect -940 2480 -720 2500
rect -940 2440 -920 2480
rect -740 2440 -720 2480
rect -940 2400 -720 2440
rect -660 2480 -440 2500
rect -660 2440 -640 2480
rect -460 2440 -440 2480
rect -660 2400 -440 2440
rect -380 2480 -160 2500
rect -380 2440 -360 2480
rect -180 2440 -160 2480
rect -380 2400 -160 2440
rect -1220 360 -1000 400
rect -1220 320 -1200 360
rect -1020 320 -1000 360
rect -1220 300 -1000 320
rect -940 360 -720 400
rect -940 320 -920 360
rect -740 320 -720 360
rect -940 300 -720 320
rect -660 360 -440 400
rect -660 320 -640 360
rect -460 320 -440 360
rect -660 300 -440 320
rect -380 360 -160 400
rect -380 320 -360 360
rect -180 320 -160 360
rect -380 300 -160 320
<< polycont >>
rect -1200 2440 -1020 2480
rect -920 2440 -740 2480
rect -640 2440 -460 2480
rect -360 2440 -180 2480
rect -1200 320 -1020 360
rect -920 320 -740 360
rect -640 320 -460 360
rect -360 320 -180 360
<< locali >>
rect -1220 2440 -1200 2480
rect -1020 2440 -1000 2480
rect -940 2440 -920 2480
rect -740 2440 -720 2480
rect -660 2440 -640 2480
rect -460 2440 -440 2480
rect -380 2440 -360 2480
rect -180 2440 -160 2480
rect -1270 2380 -1230 2405
rect -1270 420 -1265 2380
rect -1231 420 -1230 2380
rect -1270 395 -1230 420
rect -990 2380 -950 2405
rect -990 420 -985 2380
rect -951 420 -950 2380
rect -990 395 -950 420
rect -710 2380 -670 2405
rect -710 420 -705 2380
rect -671 420 -670 2380
rect -710 395 -670 420
rect -430 2380 -390 2405
rect -430 420 -425 2380
rect -391 420 -390 2380
rect -430 395 -390 420
rect -150 2380 -110 2405
rect -150 420 -145 2380
rect -111 420 -110 2380
rect -150 395 -110 420
rect -1220 320 -1200 360
rect -1020 320 -1000 360
rect -940 320 -920 360
rect -740 320 -720 360
rect -660 320 -640 360
rect -460 320 -440 360
rect -380 320 -360 360
rect -180 320 -160 360
<< viali >>
rect -1200 2440 -1020 2480
rect -920 2440 -740 2480
rect -640 2440 -460 2480
rect -360 2440 -180 2480
rect -1265 420 -1231 2380
rect -985 420 -951 2380
rect -705 420 -671 2380
rect -425 420 -391 2380
rect -145 420 -111 2380
rect -1200 320 -1020 360
rect -920 320 -740 360
rect -640 320 -460 360
rect -360 320 -180 360
<< metal1 >>
rect -1210 2480 -1010 2490
rect -930 2480 -730 2490
rect -650 2480 -450 2490
rect -370 2480 -170 2490
rect -1220 2440 -1200 2480
rect -1020 2440 -1000 2480
rect -940 2440 -920 2480
rect -740 2440 -720 2480
rect -660 2440 -640 2480
rect -460 2440 -440 2480
rect -380 2440 -360 2480
rect -180 2440 -160 2480
rect -1210 2430 -1010 2440
rect -930 2430 -730 2440
rect -650 2430 -450 2440
rect -370 2430 -170 2440
rect -1275 2380 -1225 2400
rect -1275 420 -1265 2380
rect -1231 420 -1225 2380
rect -1275 400 -1225 420
rect -995 2380 -945 2400
rect -995 420 -985 2380
rect -951 420 -945 2380
rect -995 400 -945 420
rect -715 2380 -665 2400
rect -715 420 -705 2380
rect -671 420 -665 2380
rect -715 400 -665 420
rect -435 2380 -385 2400
rect -435 420 -425 2380
rect -391 420 -385 2380
rect -435 400 -385 420
rect -155 2380 -105 2400
rect -155 420 -145 2380
rect -111 420 -105 2380
rect -155 400 -105 420
rect -1210 360 -1010 370
rect -930 360 -730 370
rect -650 360 -450 370
rect -370 360 -170 370
rect -1220 320 -1200 360
rect -1020 320 -1000 360
rect -940 320 -920 360
rect -740 320 -720 360
rect -660 320 -640 360
rect -460 320 -440 360
rect -380 320 -360 360
rect -180 320 -160 360
rect -1210 310 -1010 320
rect -930 310 -730 320
rect -650 310 -450 320
rect -370 310 -170 320
use sky130_fd_pr__nfet_01v8_TCXCTP  sky130_fd_pr__nfet_01v8_TCXCTP_0
timestamp 1728490836
transform 1 0 1095 0 1 1400
box -683 -1210 683 1210
<< end >>
