magic
tech sky130A
timestamp 1732727299
<< nwell >>
rect -500 -1000 600 300
<< pmos >>
rect -200 0 400 100
rect -200 -200 400 -100
rect -200 -400 400 -300
rect -200 -600 400 -500
rect -200 -800 400 -700
<< pdiff >>
rect -200 180 400 200
rect -200 120 -180 180
rect 380 120 400 180
rect -200 100 400 120
rect -200 -20 400 0
rect -200 -80 -180 -20
rect 380 -80 400 -20
rect -200 -100 400 -80
rect -200 -220 400 -200
rect -200 -280 -180 -220
rect 380 -280 400 -220
rect -200 -300 400 -280
rect -200 -420 400 -400
rect -200 -480 -180 -420
rect 380 -480 400 -420
rect -200 -500 400 -480
rect -200 -620 400 -600
rect -200 -680 -180 -620
rect 380 -680 400 -620
rect -200 -700 400 -680
rect -200 -820 400 -800
rect -200 -880 -180 -820
rect 380 -880 400 -820
rect -200 -900 400 -880
<< pdiffc >>
rect -180 120 380 180
rect -180 -80 380 -20
rect -180 -280 380 -220
rect -180 -480 380 -420
rect -180 -680 380 -620
rect -180 -880 380 -820
<< poly >>
rect -450 80 -200 100
rect -450 -780 -430 80
rect -370 0 -200 80
rect 400 0 500 100
rect -370 -100 -300 0
rect -370 -200 -200 -100
rect 400 -200 500 -100
rect -370 -300 -300 -200
rect -370 -400 -200 -300
rect 400 -400 500 -300
rect -370 -500 -350 -400
rect -370 -600 -200 -500
rect 400 -600 500 -500
rect -370 -700 -300 -600
rect -370 -780 -200 -700
rect -450 -800 -200 -780
rect 400 -800 500 -700
<< polycont >>
rect -430 -780 -370 80
<< locali >>
rect -300 180 400 200
rect -300 120 -180 180
rect 380 120 400 180
rect -300 100 400 120
rect -450 80 -350 100
rect -450 -780 -430 80
rect -370 -780 -350 80
rect -300 -200 -250 100
rect -200 -20 500 0
rect -200 -80 -180 -20
rect 380 -80 500 -20
rect -200 -100 500 -80
rect -300 -220 400 -200
rect -300 -280 -180 -220
rect 380 -280 400 -220
rect -300 -300 400 -280
rect -300 -600 -250 -300
rect 450 -400 500 -100
rect -200 -420 500 -400
rect -200 -480 -180 -420
rect 380 -480 500 -420
rect -200 -500 500 -480
rect -300 -620 400 -600
rect -300 -680 -180 -620
rect 380 -680 400 -620
rect -300 -700 400 -680
rect -450 -800 -350 -780
rect 450 -800 500 -500
rect -200 -820 500 -800
rect -200 -880 -180 -820
rect 380 -880 500 -820
rect -200 -900 500 -880
<< labels >>
flabel pdiffc 90 150 90 150 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont -400 -350 -400 -350 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel pdiffc 110 -850 110 -850 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell -400 210 -400 210 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
