magic
tech sky130A
magscale 1 2
timestamp 1732738914
<< nmos >>
rect -100 -269 100 331
<< ndiff >>
rect -158 319 -100 331
rect -158 -257 -146 319
rect -112 -257 -100 319
rect -158 -269 -100 -257
rect 100 319 158 331
rect 100 -257 112 319
rect 146 -257 158 319
rect 100 -269 158 -257
<< ndiffc >>
rect -146 -257 -112 319
rect 112 -257 146 319
<< poly >>
rect -100 331 100 357
rect -100 -307 100 -269
rect -100 -341 -84 -307
rect 84 -341 100 -307
rect -100 -357 100 -341
<< polycont >>
rect -84 -341 84 -307
<< locali >>
rect -146 319 -112 335
rect -146 -273 -112 -257
rect 112 319 146 335
rect 112 -273 146 -257
rect -100 -341 -84 -307
rect 84 -341 100 -307
<< viali >>
rect -146 -257 -112 319
rect 112 -257 146 319
rect -84 -341 84 -307
<< metal1 >>
rect -152 319 -106 331
rect -152 -257 -146 319
rect -112 -257 -106 319
rect -152 -269 -106 -257
rect 106 319 152 331
rect 106 -257 112 319
rect 146 -257 152 319
rect 106 -269 152 -257
rect -96 -307 96 -301
rect -96 -341 -84 -307
rect 84 -341 96 -307
rect -96 -347 96 -341
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_QX7BC3 parameters
<< end >>
