magic
tech sky130A
magscale 1 2
timestamp 1732120016
<< pwell >>
rect -5600 5066 18400 6800
rect -5600 2866 162 5066
rect 4762 2866 18400 5066
rect -5600 -1200 18400 2866
<< psubdiff >>
rect -5600 6700 18400 6800
rect -5600 6500 -5200 6700
rect 18200 6500 18400 6700
rect -5600 6400 18400 6500
rect -5600 -700 -5500 6400
rect -5300 -700 -5200 6400
rect -5600 -800 -5200 -700
rect 18000 6300 18400 6400
rect 18000 -800 18100 6300
rect 18300 -800 18400 6300
rect -5600 -900 18400 -800
rect -5600 -1100 -5400 -900
rect 17800 -1100 18400 -900
rect -5600 -1200 18400 -1100
<< psubdiffcont >>
rect -5200 6500 18200 6700
rect -5500 -700 -5300 6400
rect 18100 -800 18300 6300
rect -5400 -1100 17800 -900
<< locali >>
rect -5600 6700 18400 6800
rect -5600 6500 -5200 6700
rect 18200 6500 18400 6700
rect -5600 6400 18400 6500
rect -5600 -700 -5500 6400
rect -5300 4200 -2600 6400
rect 18000 6300 18400 6400
rect -5300 -700 -5200 4200
rect -680 2980 -280 3000
rect -680 2780 -660 2980
rect -680 2550 -280 2780
rect -3070 2440 130 2550
rect -5600 -800 -5200 -700
rect -4640 -800 -3500 -300
rect -400 -800 600 -400
rect 5400 -500 17700 -300
rect 5400 -600 11400 -500
rect 11700 -600 17700 -500
rect 5400 -800 17700 -600
rect 18000 -800 18100 6300
rect 18300 -800 18400 6300
rect -5600 -900 18400 -800
rect -5600 -1100 -5400 -900
rect 17800 -1100 18400 -900
rect -5600 -1200 18400 -1100
<< viali >>
rect -5200 6500 18200 6700
rect -5500 -700 -5300 6400
rect -900 5600 0 5800
rect -2200 5400 -1400 5600
rect 1462 4916 3262 5016
rect 900 4740 1620 4780
rect 3060 4740 3940 4780
rect -4530 3690 -3650 3950
rect 1340 3230 1460 3290
rect 3590 3230 3730 3290
rect -2240 2920 -1540 3160
rect -660 2780 -260 2980
rect 1300 2600 1500 2700
rect 3610 2630 3730 2690
rect -3310 1910 -3210 2180
rect -468 410 -434 2386
rect -210 410 -176 2386
rect 4930 1720 5030 1980
rect -10 820 70 910
rect 4940 860 5020 1020
rect -406 326 -238 360
rect -50 120 70 160
rect 3090 -220 3400 -180
rect -1340 -460 -1040 -360
rect 11400 -600 11700 -500
rect 18100 -800 18300 6300
rect -5400 -1100 17800 -900
<< metal1 >>
rect -5600 6700 18400 6800
rect -5600 6500 -5200 6700
rect 18200 6500 18400 6700
rect -5600 6400 18400 6500
rect -5600 -700 -5500 6400
rect -5300 4200 -2600 6400
rect 18000 6300 18400 6400
rect -2500 5800 4500 6300
rect -2500 5600 -900 5800
rect 0 5600 4500 5800
rect -2500 5400 -2200 5600
rect -1400 5400 4500 5600
rect -2500 5300 -1200 5400
rect 640 5016 4500 5400
rect 212 4916 1462 5016
rect 3262 4916 4712 5016
rect -5300 -700 -5200 4200
rect -4640 3950 -2540 4030
rect -4640 3690 -4530 3950
rect -3650 3690 -2540 3950
rect -4640 3660 -2540 3690
rect -3360 3260 -2550 3660
rect -3360 3160 -1280 3260
rect -3360 2920 -2240 3160
rect -1540 2920 -1280 3160
rect 212 3066 312 4916
rect 640 4780 4500 4916
rect 640 4740 900 4780
rect 1620 4740 3060 4780
rect 3940 4740 4500 4780
rect 640 4720 4500 4740
rect 1320 3290 1480 3310
rect 1320 3230 1340 3290
rect 1460 3230 1480 3290
rect 1320 3210 1480 3230
rect 3570 3290 3770 3310
rect 3570 3230 3590 3290
rect 3730 3230 3770 3290
rect 3570 3220 3770 3230
rect 4612 3066 4712 4916
rect -3360 2820 -1280 2920
rect -680 2980 -240 3000
rect -3360 2180 -3170 2820
rect -680 2780 -660 2980
rect -260 2780 -240 2980
rect 212 2966 4712 3066
rect -680 2760 -240 2780
rect 1280 2700 1520 2720
rect 1280 2600 1300 2700
rect 1500 2600 1520 2700
rect 3590 2690 3750 2710
rect 3590 2630 3610 2690
rect 3730 2630 3750 2690
rect 3590 2610 3750 2630
rect 1280 2580 1520 2600
rect -3360 1910 -3310 2180
rect -3210 1910 -3170 2180
rect -3360 1730 -3170 1910
rect 4910 1980 5050 1990
rect 4910 1720 4930 1980
rect 5030 1720 5050 1980
rect 4910 1710 5050 1720
rect 4870 1020 5110 1100
rect -70 910 90 920
rect -70 820 -10 910
rect 70 820 90 910
rect -176 410 -100 440
rect -420 300 -410 370
rect -230 300 -220 370
rect -420 290 -220 300
rect -140 260 -100 410
rect -210 230 -100 260
rect -5600 -800 -5200 -700
rect -4640 -800 -3500 -300
rect -1380 -360 -980 -340
rect -1380 -460 -1340 -360
rect -1040 -460 -980 -360
rect -210 -400 -160 230
rect -70 160 90 820
rect 4870 860 4940 1020
rect 5020 860 5110 1020
rect 120 540 200 550
rect 120 360 130 540
rect 120 350 200 360
rect -70 120 -50 160
rect 70 120 90 160
rect -70 110 90 120
rect 370 -400 480 322
rect 4870 -150 5110 860
rect 3030 -180 5110 -150
rect 3030 -220 3090 -180
rect 3400 -220 5110 -180
rect 3030 -230 5110 -220
rect -1380 -480 -980 -460
rect -1340 -640 -1040 -480
rect -400 -800 600 -400
rect 5400 -500 17700 -300
rect 5400 -600 11400 -500
rect 11700 -600 17700 -500
rect 5400 -800 17700 -600
rect 18000 -800 18100 6300
rect 18300 -800 18400 6300
rect -5600 -900 18400 -800
rect -5600 -1100 -5400 -900
rect 17800 -1100 18400 -900
rect -5600 -1200 18400 -1100
<< via1 >>
rect 1340 3230 1460 3290
rect 3590 3230 3730 3290
rect 1300 2600 1500 2700
rect 3610 2630 3730 2690
rect 4930 1720 5030 1980
rect -410 360 -230 370
rect -410 326 -406 360
rect -406 326 -238 360
rect -238 326 -230 360
rect -410 300 -230 326
rect 130 360 200 540
rect 11400 -600 11700 -500
<< metal2 >>
rect 1300 3290 1500 3310
rect 1300 3230 1340 3290
rect 1460 3230 1500 3290
rect 1300 2720 1500 3230
rect 3570 3290 3770 3310
rect 3570 3230 3590 3290
rect 3730 3230 3770 3290
rect 3570 3220 3770 3230
rect 1280 2700 1520 2720
rect 1280 2600 1300 2700
rect 1500 2600 1520 2700
rect 3590 2690 3750 3220
rect 3590 2630 3610 2690
rect 3730 2630 3750 2690
rect 3590 2610 3750 2630
rect 1280 2580 1520 2600
rect 4910 1980 5050 1990
rect 4910 1720 4930 1980
rect 5030 1720 5050 1980
rect 4910 1710 5050 1720
rect 110 540 210 550
rect 110 380 130 540
rect -420 370 130 380
rect -420 300 -410 370
rect -230 360 130 370
rect 200 360 210 540
rect -230 300 210 360
rect -420 290 -220 300
rect 11300 -500 11800 -400
rect 11300 -600 11400 -500
rect 11700 -600 11800 -500
rect 11300 -700 11800 -600
<< via2 >>
rect 4930 1720 5030 1980
rect 11400 -600 11700 -500
<< metal3 >>
rect 4910 1980 5050 1990
rect 4910 1720 4930 1980
rect 5030 1720 5050 1980
rect 4910 1710 5050 1720
rect 11300 -500 11800 -400
rect 11300 -600 11400 -500
rect 11700 -600 11800 -500
rect 11300 -700 11800 -600
<< via3 >>
rect 4930 1720 5030 1980
rect 11400 -600 11700 -500
<< metal4 >>
rect 10800 3000 12000 3800
rect 4900 1980 5700 2000
rect 4900 1720 4930 1980
rect 5030 1720 5700 1980
rect 4900 1700 5700 1720
rect 11300 -200 11800 -100
rect 11500 -400 11600 -200
rect 11300 -500 11800 -400
rect 11300 -600 11400 -500
rect 11700 -600 11800 -500
rect 11300 -700 11800 -600
use diff_pair_n  diff_pair_n_0
timestamp 1731518228
transform 1 0 1680 0 1 1460
box -1800 -1000 3450 1400
use diff_pair_p  diff_pair_p_0
timestamp 1731631080
transform -1 0 3362 0 -1 3866
box -1400 -1200 3200 1000
use n70x1  n70x1_0
timestamp 1731632322
transform 1 0 -1960 0 1 1500
box -1800 -2200 1800 1200
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1731631080
transform 0 1 8440 -1 0 2986
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_1
timestamp 1731631080
transform 0 1 14640 -1 0 2986
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_7JY9FK  sky130_fd_pr__nfet_01v8_7JY9FK_0
timestamp 1731632322
transform -1 0 -322 0 1 1367
box -158 -1057 158 1057
use sky130_fd_pr__nfet_01v8_QX7BC3  sky130_fd_pr__nfet_01v8_QX7BC3_0
timestamp 1732120016
transform 0 1 501 -1 0 428
box -158 -357 158 357
use sky130_fd_pr__res_xhigh_po_0p35_BB2ZH9  sky130_fd_pr__res_xhigh_po_0p35_BB2ZH9_0
timestamp 1732120016
transform 0 1 1670 -1 0 -47
box -201 -1796 201 1796
use sky130_fd_pr__res_xhigh_po_5p73_7D764L  sky130_fd_pr__res_xhigh_po_5p73_7D764L_0
timestamp 1731631080
transform 1 0 -467 0 1 4296
box -573 -1616 573 1616
use sky130_fd_pr__res_xhigh_po_5p73_F3YNPN  sky130_fd_pr__res_xhigh_po_5p73_F3YNPN_0
timestamp 1731631080
transform 1 0 -1837 0 1 4266
box -573 -1416 573 1416
use sky130_fd_pr__res_xhigh_po_5p73_G7VZ5E  sky130_fd_pr__res_xhigh_po_5p73_G7VZ5E_0
timestamp 1731631080
transform 1 0 -4067 0 1 1716
box -573 -2416 573 2416
<< labels >>
flabel metal1 1600 5700 1600 5700 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel via1 3660 2660 3660 2660 0 FreeSans 1600 0 0 0 Voutp
port 2 nsew
flabel via1 1320 2660 1320 2660 0 FreeSans 1600 0 0 0 Voutn
port 1 nsew
flabel metal1 5020 460 5020 460 0 FreeSans 1600 0 0 0 Vg3
flabel via1 -280 340 -280 340 0 FreeSans 1600 0 0 0 Vref
port 4 nsew
flabel locali -460 2520 -460 2520 0 FreeSans 1600 0 0 0 Vg2
flabel metal1 -2920 3380 -2920 3380 0 FreeSans 1600 0 0 0 Vg
flabel viali -3100 6600 -3100 6600 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel metal1 -1200 -560 -1200 -560 0 FreeSans 1600 0 0 0 Vin
port 3 nsew
<< end >>
