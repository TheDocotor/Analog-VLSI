magic
tech sky130A
magscale 1 2
timestamp 1726675666
<< pwell >>
rect -2306 -98 -908 2292
<< nmos >>
rect -2080 104 -1130 2076
<< ndiff >>
rect -2152 2014 -2080 2076
rect -2152 168 -2134 2014
rect -2098 168 -2080 2014
rect -2152 104 -2080 168
rect -1130 1978 -1050 2076
rect -1130 154 -1106 1978
rect -1072 154 -1050 1978
rect -1130 104 -1050 154
<< ndiffc >>
rect -2134 168 -2098 2014
rect -1106 154 -1072 1978
<< psubdiff >>
rect -2266 2202 -2152 2248
rect -1042 2202 -946 2248
rect -2266 2140 -2222 2202
rect -980 2130 -946 2202
rect -2266 -26 -2222 30
rect -980 -26 -946 58
rect -2266 -60 -2136 -26
rect -1042 -60 -946 -26
<< psubdiffcont >>
rect -2152 2202 -1042 2248
rect -2266 30 -2222 2140
rect -980 58 -946 2130
rect -2136 -60 -1042 -26
<< poly >>
rect -2080 2148 -1130 2166
rect -2080 2114 -2044 2148
rect -1154 2114 -1130 2148
rect -2080 2076 -1130 2114
rect -2080 66 -1130 104
rect -2080 32 -2044 66
rect -1154 32 -1130 66
rect -2080 10 -1130 32
<< polycont >>
rect -2044 2114 -1154 2148
rect -2044 32 -1154 66
<< locali >>
rect -2262 2244 -2152 2248
rect -2266 2202 -2152 2244
rect -1042 2202 -946 2248
rect -2266 2140 -2222 2202
rect -2080 2114 -2044 2148
rect -1154 2114 -1130 2148
rect -980 2130 -946 2202
rect -2134 2014 -2098 2076
rect -2134 98 -2098 168
rect -1106 1978 -1070 2074
rect -1072 154 -1070 1978
rect -1106 104 -1070 154
rect -2080 32 -2044 66
rect -1154 32 -1130 66
rect -2266 -26 -2222 30
rect -980 -26 -946 58
rect -2266 -60 -2136 -26
rect -1042 -60 -946 -26
<< viali >>
rect -2044 2114 -1154 2148
rect -2134 168 -2098 2014
rect -1106 154 -1072 1978
rect -2044 32 -1154 66
<< metal1 >>
rect -2072 2148 -1140 2156
rect -2072 2114 -2044 2148
rect -1154 2114 -1140 2148
rect -2072 2100 -1140 2114
rect -2142 2014 -2090 2076
rect -2142 168 -2134 2014
rect -2098 168 -2090 2014
rect -2142 104 -2090 168
rect -1116 1978 -1060 2076
rect -1116 154 -1106 1978
rect -1072 154 -1060 1978
rect -1116 104 -1060 154
rect -2064 66 -1140 76
rect -2064 32 -2044 66
rect -1154 32 -1140 66
rect -2064 26 -1140 32
use sky130_fd_pr__nfet_01v8_TSEK3K  sky130_fd_pr__nfet_01v8_TSEK3K_0
timestamp 1726675666
transform 1 0 1569 0 1 1751
box -696 -1210 696 1210
<< end >>
