magic
tech sky130A
magscale 1 2
timestamp 1729279979
<< xpolycontact >>
rect -69 329 69 761
rect -69 -761 69 -329
<< xpolyres >>
rect -69 -329 69 329
<< viali >>
rect -53 346 53 743
rect -53 -743 53 -346
<< metal1 >>
rect -59 743 59 755
rect -59 346 -53 743
rect 53 346 59 743
rect -59 334 59 346
rect -59 -346 59 -334
rect -59 -743 -53 -346
rect 53 -743 59 -346
rect -59 -755 59 -743
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.69 l 3.45 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 10.545k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_0p69_2LTKQM parameters
<< end >>
