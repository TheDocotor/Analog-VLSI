magic
tech sky130A
timestamp 1732726409
<< nwell >>
rect -500 -600 500 300
<< pmos >>
rect -200 0 300 100
rect -200 -200 300 -100
rect -200 -400 300 -300
<< pdiff >>
rect -200 180 300 200
rect -200 120 -180 180
rect 280 120 300 180
rect -200 100 300 120
rect -200 -20 300 0
rect -200 -80 -180 -20
rect 280 -80 300 -20
rect -200 -100 300 -80
rect -200 -220 300 -200
rect -200 -280 -180 -220
rect 280 -280 300 -220
rect -200 -300 300 -280
rect -200 -420 300 -400
rect -200 -480 -180 -420
rect 280 -480 300 -420
rect -200 -500 300 -480
<< pdiffc >>
rect -180 120 280 180
rect -180 -80 280 -20
rect -180 -280 280 -220
rect -180 -480 280 -420
<< poly >>
rect -450 80 -200 100
rect -450 -380 -430 80
rect -370 0 -200 80
rect 300 0 400 100
rect -370 -100 -300 0
rect -370 -200 -200 -100
rect 300 -200 400 -100
rect -370 -300 -300 -200
rect -370 -380 -200 -300
rect -450 -400 -200 -380
rect 300 -400 400 -300
<< polycont >>
rect -430 -380 -370 80
<< locali >>
rect -300 180 300 200
rect -300 120 -180 180
rect 280 120 300 180
rect -300 100 300 120
rect -450 80 -350 100
rect -450 -380 -430 80
rect -370 -380 -350 80
rect -300 -200 -250 100
rect -200 -20 400 0
rect -200 -80 -180 -20
rect 280 -80 400 -20
rect -200 -100 400 -80
rect -300 -220 300 -200
rect -300 -280 -180 -220
rect 280 -280 300 -220
rect -300 -300 300 -280
rect -450 -400 -350 -380
rect 350 -400 400 -100
rect -200 -420 400 -400
rect -200 -480 -180 -420
rect 280 -480 400 -420
rect -200 -500 400 -480
<< labels >>
flabel pdiffc 40 150 40 150 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont -400 -150 -400 -150 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel pdiffc 60 -450 60 -450 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell -400 210 -400 210 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
