magic
tech sky130A
magscale 1 2
timestamp 1731517860
<< nwell >>
rect -225 -1150 1875 550
<< pmos >>
rect 100 200 1700 400
rect 100 -100 1700 100
rect 100 -400 1700 -200
rect 100 -700 1700 -500
rect 100 -1000 1700 -800
<< pdiff >>
rect 100 475 1700 500
rect 100 425 125 475
rect 1675 425 1700 475
rect 100 400 1700 425
rect 100 175 1700 200
rect 100 125 125 175
rect 1675 125 1700 175
rect 100 100 1700 125
rect 100 -125 1700 -100
rect 100 -175 125 -125
rect 1675 -175 1700 -125
rect 100 -200 1700 -175
rect 100 -425 1700 -400
rect 100 -475 125 -425
rect 1675 -475 1700 -425
rect 100 -500 1700 -475
rect 100 -725 1700 -700
rect 100 -775 125 -725
rect 1675 -775 1700 -725
rect 100 -800 1700 -775
rect 100 -1025 1700 -1000
rect 100 -1075 125 -1025
rect 1675 -1075 1700 -1025
rect 100 -1100 1700 -1075
<< pdiffc >>
rect 125 425 1675 475
rect 125 125 1675 175
rect 125 -175 1675 -125
rect 125 -475 1675 -425
rect 125 -775 1675 -725
rect 125 -1075 1675 -1025
<< poly >>
rect -200 375 100 400
rect -200 -975 -175 375
rect -125 200 100 375
rect 1700 200 1800 400
rect -125 100 0 200
rect -125 -100 100 100
rect 1700 -100 1800 100
rect -125 -200 0 -100
rect -125 -400 100 -200
rect 1700 -400 1800 -200
rect -125 -500 0 -400
rect -125 -700 100 -500
rect 1700 -700 1800 -500
rect -125 -800 0 -700
rect -125 -975 100 -800
rect -200 -1000 100 -975
rect 1700 -1000 1800 -800
<< polycont >>
rect -175 -975 -125 375
<< locali >>
rect -50 475 1700 500
rect -50 425 125 475
rect 1675 425 1700 475
rect -50 400 1700 425
rect -200 375 -100 400
rect -200 -975 -175 375
rect -125 -975 -100 375
rect -50 -100 50 400
rect 100 175 1850 200
rect 100 125 125 175
rect 1675 125 1850 175
rect 100 100 1850 125
rect -50 -125 1700 -100
rect -50 -175 125 -125
rect 1675 -175 1700 -125
rect -50 -200 1700 -175
rect -50 -700 50 -200
rect 1750 -400 1850 100
rect 100 -425 1850 -400
rect 100 -475 125 -425
rect 1675 -475 1850 -425
rect 100 -500 1850 -475
rect -50 -725 1700 -700
rect -50 -775 125 -725
rect 1675 -775 1700 -725
rect -50 -800 1700 -775
rect -200 -1000 -100 -975
rect 1750 -1000 1850 -500
rect 100 -1025 1850 -1000
rect 100 -1075 125 -1025
rect 1675 -1075 1850 -1025
rect 100 -1100 1850 -1075
<< labels >>
flabel pdiffc 600 450 600 450 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel pdiffc 625 -1050 625 -1050 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel polycont -150 -300 -150 -300 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel nwell -150 475 -150 475 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
