magic
tech sky130A
timestamp 1730605901
<< nmos >>
rect -250 -50 250 50
<< ndiff >>
rect -279 44 -250 50
rect -279 -44 -273 44
rect -256 -44 -250 44
rect -279 -50 -250 -44
rect 250 44 279 50
rect 250 -44 256 44
rect 273 -44 279 44
rect 250 -50 279 -44
<< ndiffc >>
rect -273 -44 -256 44
rect 256 -44 273 44
<< poly >>
rect -250 50 250 63
rect -250 -63 250 -50
<< locali >>
rect -273 44 -256 52
rect -273 -52 -256 -44
rect 256 44 273 52
rect 256 -52 273 -44
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_ZCPJ4U parameters
<< end >>
