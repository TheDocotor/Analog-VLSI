magic
tech sky130A
magscale 1 2
timestamp 1730605901
<< xpolycontact >>
rect 1911 1244 3057 1676
rect -3057 -1676 -1911 -1244
<< xpolyres >>
rect -3057 6 -669 1140
rect -573 6 1815 1140
rect 1911 6 3057 1244
rect -3057 -6 3057 6
rect -3057 -1244 -1911 -6
rect -1815 -1140 573 -6
rect 669 -1140 3057 -6
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 11.4 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 27.96k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_5p73_QHLGXT parameters
<< end >>
