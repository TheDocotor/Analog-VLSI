magic
tech sky130A
magscale 1 2
timestamp 1729280326
<< pwell >>
rect -235 -893 235 893
<< psubdiff >>
rect -199 823 -103 857
rect 103 823 199 857
rect -199 761 -165 823
rect 165 761 199 823
rect -199 -823 -165 -761
rect 165 -823 199 -761
rect -199 -857 -103 -823
rect 103 -857 199 -823
<< psubdiffcont >>
rect -103 823 103 857
rect -199 -761 -165 761
rect 165 -761 199 761
rect -103 -857 103 -823
<< xpolycontact >>
rect -69 295 69 727
rect -69 -727 69 -295
<< xpolyres >>
rect -69 -295 69 295
<< locali >>
rect -199 823 -103 857
rect 103 823 199 857
rect -199 761 -165 823
rect 165 761 199 823
rect -199 -823 -165 -761
rect 165 -823 199 -761
rect -199 -857 -103 -823
rect 103 -857 199 -823
<< viali >>
rect -53 312 53 709
rect -53 -709 53 -312
<< metal1 >>
rect -59 709 59 721
rect -59 312 -53 709
rect 53 312 59 709
rect -59 300 59 312
rect -59 -312 59 -300
rect -59 -709 -53 -312
rect 53 -709 59 -312
rect -59 -721 59 -709
<< properties >>
string FIXED_BBOX -182 -840 182 840
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.69 l 3.105 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 9.545k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_0p69_S6L29W parameters
<< end >>
