* SPICE3 file created from diff_pair_d.ext - technology: sky130A

.subckt nmos_40 D G S B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.3 as=1.5 ps=10.3 w=10 l=1.1
X1 D G S B sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.3 as=3 ps=20.6 w=10 l=1.1
X2 S G D B sky130_fd_pr__nfet_01v8 ad=3 pd=20.6 as=1.5 ps=10.3 w=10 l=1.1
X3 S G D B sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.3 as=1.5 ps=10.3 w=10 l=1.1
C0 S G 3.20505f
C1 D G 2.53191f
C2 S D 2.16384f
C3 G B 2.53805f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_2LTKQM a_n69_n761# a_n69_329# VSUBS
X0 a_n69_329# a_n69_n761# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt Rf_res sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1/a_n69_n761# sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_0/a_n69_329#
+ VSUBS sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1/a_n69_329#
Xsky130_fd_pr__res_xhigh_po_0p69_2LTKQM_0 sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1/a_n69_329#
+ sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_0/a_n69_329# VSUBS sky130_fd_pr__res_xhigh_po_0p69_2LTKQM
Xsky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1 sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1/a_n69_n761#
+ sky130_fd_pr__res_xhigh_po_0p69_2LTKQM_1/a_n69_329# VSUBS sky130_fd_pr__res_xhigh_po_0p69_2LTKQM
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_C432MY a_n69_n727# a_n69_295# VSUBS
X0 a_n69_295# a_n69_n727# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=3.11
.ends

.subckt CS_res sky130_fd_pr__res_xhigh_po_0p69_C432MY_0/a_n69_n727# sky130_fd_pr__res_xhigh_po_0p69_C432MY_0/a_n69_295#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_0p69_C432MY_0 sky130_fd_pr__res_xhigh_po_0p69_C432MY_0/a_n69_n727#
+ sky130_fd_pr__res_xhigh_po_0p69_C432MY_0/a_n69_295# VSUBS sky130_fd_pr__res_xhigh_po_0p69_C432MY
.ends

.subckt if_res a_n400_0# a_n400_2334# VSUBS
X0 a_n400_2334# a_n400_0# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=9.67
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_LZXZX3 a_n69_674# a_n69_n1106# VSUBS
X0 a_n69_674# a_n69_n1106# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=6.9
.ends

.subckt Vdd_res sky130_fd_pr__res_xhigh_po_0p69_LZXZX3_0/a_n69_n1106# VSUBS sky130_fd_pr__res_xhigh_po_0p69_LZXZX3_0/a_n69_674#
Xsky130_fd_pr__res_xhigh_po_0p69_LZXZX3_0 sky130_fd_pr__res_xhigh_po_0p69_LZXZX3_0/a_n69_674#
+ sky130_fd_pr__res_xhigh_po_0p69_LZXZX3_0/a_n69_n1106# VSUBS sky130_fd_pr__res_xhigh_po_0p69_LZXZX3
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_P8UVGE a_n69_122# a_n69_n554# VSUBS
X0 a_n69_122# a_n69_n554# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=1.38
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV a_n69_n761# a_n69_329# VSUBS
X0 a_n69_329# a_n69_n761# VSUBS sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt LOp_resistor sky130_fd_pr__res_xhigh_po_0p69_P8UVGE_0/a_n69_122# sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0/a_n69_329#
+ sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0/a_n69_n761# VSUBS
Xsky130_fd_pr__res_xhigh_po_0p69_P8UVGE_0 sky130_fd_pr__res_xhigh_po_0p69_P8UVGE_0/a_n69_122#
+ sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0/a_n69_329# VSUBS sky130_fd_pr__res_xhigh_po_0p69_P8UVGE
Xsky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0 sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0/a_n69_n761#
+ sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV_0/a_n69_329# VSUBS sky130_fd_pr__res_xhigh_po_0p69_Z9GMGV
.ends

.subckt Gilbert nmos_40_1/G nmos_40_1/D nmos_40_0/S nmos_40_0/G nmos_40_1/S VSUBS
Xnmos_40_0 nmos_40_1/D nmos_40_0/G nmos_40_0/S VSUBS nmos_40
Xnmos_40_1 nmos_40_1/D nmos_40_1/G nmos_40_1/S VSUBS nmos_40
C0 nmos_40_1/G VSUBS 2.53805f
C1 nmos_40_0/G VSUBS 2.53805f
.ends

.subckt diff_pair_d VDD VSS LOn LOp RFn RFp IFp IFn
Xnmos_40_2 VSS VSS Vamp VSUBS nmos_40
XRf_res_0 VSS VDD VSUBS RFp Rf_res
XCS_res_0 VSS VDD VSUBS CS_res
XRf_res_1 VSS VDD VSUBS RFn Rf_res
Xif_res_1 IFn VDD VSUBS if_res
Xif_res_0 VDD IFp VSUBS if_res
XVdd_res_0 VDD VSUBS IF++ Vdd_res
XVdd_res_1 VDD VSUBS IF-- Vdd_res
XLOp_resistor_0 VDD LOn VSS VSUBS LOp_resistor
XLOp_resistor_1 VDD LOp VSS VSUBS LOp_resistor
XGilbert_0 LOp Vmid IF-- LOn IF++ VSUBS Gilbert
XGilbert_1 LOn Vmid2 IF-- LOp IF++ VSUBS Gilbert
XGilbert_2 RFp VSS Vmid2 RFn Vmid VSUBS Gilbert
XGilbert_3 IF-- Vamp IFn IF++ IFp VSUBS Gilbert
Xnmos_40_0 VSS VSS VSS VSUBS nmos_40
Xnmos_40_1 VSS VSS VSS VSUBS nmos_40
C0 LOn LOp 3.089737f
C1 VSS RFn 2.161304f
C2 RFn RFp 2.146045f
C3 VSS RFp 2.190594f
C4 LOn VDD 4.22694f
C5 IF++ IF-- 5.905244f
C6 VSS VDD 4.840173f
C7 Vamp VSUBS 3.065262f
C8 IF-- VSUBS 7.894908f
C9 IFn VSUBS 2.019003f
C10 IF++ VSUBS 6.959948f
C11 RFn VSUBS 3.85366f
C12 LOp VSUBS 7.268859f
C13 LOn VSUBS 2.985119f
C14 VSS VSUBS 78.11744f
C15 VDD VSUBS 21.496222f
C16 RFp VSUBS 4.197855f
.ends

