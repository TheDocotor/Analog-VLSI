magic
tech sky130A
timestamp 1730605901
<< nwell >>
rect -684 -131 684 131
<< pmos >>
rect -637 -100 -587 100
rect -501 -100 -451 100
rect -365 -100 -315 100
rect -229 -100 -179 100
rect -93 -100 -43 100
rect 43 -100 93 100
rect 179 -100 229 100
rect 315 -100 365 100
rect 451 -100 501 100
rect 587 -100 637 100
<< pdiff >>
rect -666 94 -637 100
rect -666 -94 -660 94
rect -643 -94 -637 94
rect -666 -100 -637 -94
rect -587 94 -558 100
rect -587 -94 -581 94
rect -564 -94 -558 94
rect -587 -100 -558 -94
rect -530 94 -501 100
rect -530 -94 -524 94
rect -507 -94 -501 94
rect -530 -100 -501 -94
rect -451 94 -422 100
rect -451 -94 -445 94
rect -428 -94 -422 94
rect -451 -100 -422 -94
rect -394 94 -365 100
rect -394 -94 -388 94
rect -371 -94 -365 94
rect -394 -100 -365 -94
rect -315 94 -286 100
rect -315 -94 -309 94
rect -292 -94 -286 94
rect -315 -100 -286 -94
rect -258 94 -229 100
rect -258 -94 -252 94
rect -235 -94 -229 94
rect -258 -100 -229 -94
rect -179 94 -150 100
rect -179 -94 -173 94
rect -156 -94 -150 94
rect -179 -100 -150 -94
rect -122 94 -93 100
rect -122 -94 -116 94
rect -99 -94 -93 94
rect -122 -100 -93 -94
rect -43 94 -14 100
rect -43 -94 -37 94
rect -20 -94 -14 94
rect -43 -100 -14 -94
rect 14 94 43 100
rect 14 -94 20 94
rect 37 -94 43 94
rect 14 -100 43 -94
rect 93 94 122 100
rect 93 -94 99 94
rect 116 -94 122 94
rect 93 -100 122 -94
rect 150 94 179 100
rect 150 -94 156 94
rect 173 -94 179 94
rect 150 -100 179 -94
rect 229 94 258 100
rect 229 -94 235 94
rect 252 -94 258 94
rect 229 -100 258 -94
rect 286 94 315 100
rect 286 -94 292 94
rect 309 -94 315 94
rect 286 -100 315 -94
rect 365 94 394 100
rect 365 -94 371 94
rect 388 -94 394 94
rect 365 -100 394 -94
rect 422 94 451 100
rect 422 -94 428 94
rect 445 -94 451 94
rect 422 -100 451 -94
rect 501 94 530 100
rect 501 -94 507 94
rect 524 -94 530 94
rect 501 -100 530 -94
rect 558 94 587 100
rect 558 -94 564 94
rect 581 -94 587 94
rect 558 -100 587 -94
rect 637 94 666 100
rect 637 -94 643 94
rect 660 -94 666 94
rect 637 -100 666 -94
<< pdiffc >>
rect -660 -94 -643 94
rect -581 -94 -564 94
rect -524 -94 -507 94
rect -445 -94 -428 94
rect -388 -94 -371 94
rect -309 -94 -292 94
rect -252 -94 -235 94
rect -173 -94 -156 94
rect -116 -94 -99 94
rect -37 -94 -20 94
rect 20 -94 37 94
rect 99 -94 116 94
rect 156 -94 173 94
rect 235 -94 252 94
rect 292 -94 309 94
rect 371 -94 388 94
rect 428 -94 445 94
rect 507 -94 524 94
rect 564 -94 581 94
rect 643 -94 660 94
<< poly >>
rect -637 100 -587 113
rect -501 100 -451 113
rect -365 100 -315 113
rect -229 100 -179 113
rect -93 100 -43 113
rect 43 100 93 113
rect 179 100 229 113
rect 315 100 365 113
rect 451 100 501 113
rect 587 100 637 113
rect -637 -113 -587 -100
rect -501 -113 -451 -100
rect -365 -113 -315 -100
rect -229 -113 -179 -100
rect -93 -113 -43 -100
rect 43 -113 93 -100
rect 179 -113 229 -100
rect 315 -113 365 -100
rect 451 -113 501 -100
rect 587 -113 637 -100
<< locali >>
rect -660 94 -643 102
rect -660 -102 -643 -94
rect -581 94 -564 102
rect -581 -102 -564 -94
rect -524 94 -507 102
rect -524 -102 -507 -94
rect -445 94 -428 102
rect -445 -102 -428 -94
rect -388 94 -371 102
rect -388 -102 -371 -94
rect -309 94 -292 102
rect -309 -102 -292 -94
rect -252 94 -235 102
rect -252 -102 -235 -94
rect -173 94 -156 102
rect -173 -102 -156 -94
rect -116 94 -99 102
rect -116 -102 -99 -94
rect -37 94 -20 102
rect -37 -102 -20 -94
rect 20 94 37 102
rect 20 -102 37 -94
rect 99 94 116 102
rect 99 -102 116 -94
rect 156 94 173 102
rect 156 -102 173 -94
rect 235 94 252 102
rect 235 -102 252 -94
rect 292 94 309 102
rect 292 -102 309 -94
rect 371 94 388 102
rect 371 -102 388 -94
rect 428 94 445 102
rect 428 -102 445 -94
rect 507 94 524 102
rect 507 -102 524 -94
rect 564 94 581 102
rect 564 -102 581 -94
rect 643 94 660 102
rect 643 -102 660 -94
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l .5 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_01v8_URPVEG parameters
<< end >>
