magic
tech sky130A
magscale 1 2
timestamp 1732122809
<< nmos >>
rect -800 -531 800 469
<< ndiff >>
rect -858 457 -800 469
rect -858 -519 -846 457
rect -812 -519 -800 457
rect -858 -531 -800 -519
rect 800 457 858 469
rect 800 -519 812 457
rect 846 -519 858 457
rect 800 -531 858 -519
<< ndiffc >>
rect -846 -519 -812 457
rect 812 -519 846 457
<< poly >>
rect -800 541 800 557
rect -800 507 -784 541
rect 784 507 800 541
rect -800 469 800 507
rect -800 -557 800 -531
<< polycont >>
rect -784 507 784 541
<< locali >>
rect -800 507 -784 541
rect 784 507 800 541
rect -846 457 -812 473
rect -846 -535 -812 -519
rect 812 457 846 473
rect 812 -535 846 -519
<< viali >>
rect -784 507 784 541
rect -846 -519 -812 457
rect 812 -519 846 457
<< metal1 >>
rect -796 541 796 547
rect -796 507 -784 541
rect 784 507 796 541
rect -796 501 796 507
rect -852 457 -806 469
rect -852 -519 -846 457
rect -812 -519 -806 457
rect -852 -531 -806 -519
rect 806 457 852 469
rect 806 -519 812 457
rect 846 -519 852 457
rect 806 -531 852 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_8K47H6 parameters
<< end >>
