magic
tech sky130A
magscale 1 2
timestamp 1730767210
<< pwell >>
rect -739 -8582 739 8582
<< psubdiff >>
rect -703 8512 -607 8546
rect 607 8512 703 8546
rect -703 8450 -669 8512
rect 669 8450 703 8512
rect -703 -8512 -669 -8450
rect 669 -8512 703 -8450
rect -703 -8546 -607 -8512
rect 607 -8546 703 -8512
<< psubdiffcont >>
rect -607 8512 607 8546
rect -703 -8450 -669 8450
rect 669 -8450 703 8450
rect -607 -8546 607 -8512
<< xpolycontact >>
rect -573 7984 573 8416
rect -573 -8416 573 -7984
<< xpolyres >>
rect -573 -7984 573 7984
<< locali >>
rect -703 8512 -607 8546
rect 607 8512 703 8546
rect -703 8450 -669 8512
rect 669 8450 703 8512
rect -703 -8512 -669 -8450
rect 669 -8512 703 -8450
rect -703 -8546 -607 -8512
rect 607 -8546 703 -8512
<< viali >>
rect -557 8001 557 8398
rect -557 -8398 557 -8001
<< metal1 >>
rect -569 8398 569 8404
rect -569 8001 -557 8398
rect 557 8001 569 8398
rect -569 7995 569 8001
rect -569 -8001 569 -7995
rect -569 -8398 -557 -8001
rect 557 -8398 569 -8001
rect -569 -8404 569 -8398
<< properties >>
string FIXED_BBOX -686 -8529 686 8529
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 80 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 27.988k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_5p73_X7VN8P parameters
<< end >>
