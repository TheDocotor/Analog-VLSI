** sch_path: /home/renslow/Documents/ece5120/hw02/xschem/amp_tb.sch
**.subckt amp_tb
V1 net1 GND 5.0
V2 Vin GND ac 1 sine(0 5m 1k)
x1 net1 Vout Vin GND cs_amp
R1 Vout GND 1Meg m=1
**** begin user architecture code



.option wnflag=1
.option savecurrents
.include ../mag/my_nmos.spice

.control
save all
tran 10u 2m
set color0=white
set color1=blue
plot vin, vout
ac dec 100 10 1000meg
let mag = db(vout)
plot mag
let phase = cph(vout)*180/pi
plot phase
save all
write hw1_tb.raw

.endc



** opencircuitdesign pdks install
.lib /usr/magic/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  cs_amp.sym # of pins=4
** sym_path: /home/renslow/Documents/ece5120/hw02/xschem/cs_amp.sym
** sch_path: /home/renslow/Documents/ece5120/hw02/xschem/cs_amp.sch
.subckt cs_amp VDD Vo Vin VSS
*.ipin Vin
*.ipin VDD
*.opin Vo
*.ipin VSS
x1 V_D V_gate net1 VSS my_nmos
C1 Vin V_gate 100u m=1
C2 Vo V_D 100u m=1
Vmeas net1 VSS 0
.save i(vmeas)
R1 VDD V_gate 400k m=1
R2 V_gate VSS 100k m=1
R3 VDD V_D 76.9k m=1
.ends

.GLOBAL GND
.end
