magic
tech sky130A
magscale 1 2
timestamp 1730316371
<< nwell >>
rect -2200 4400 6000 5400
<< mvnsubdiff >>
rect -2120 5180 5920 5280
rect -2120 4560 -2040 5180
rect 5840 4560 5920 5180
rect -2120 4480 5920 4560
<< locali >>
rect -2120 5180 5920 5280
rect -2120 4560 -2040 5180
rect 5840 4560 5920 5180
rect -2120 4480 5920 4560
rect 2020 420 2180 1580
<< viali >>
rect 1120 3600 1280 3640
<< metal1 >>
rect -2200 5120 6000 5640
rect -2120 4560 -2040 5120
rect 1100 4900 1300 5120
rect 1100 4560 1300 4680
rect 5840 4560 5920 5120
rect -2120 4480 5920 4560
rect 1100 3640 1300 4480
rect 1100 3600 1120 3640
rect 1280 3600 1300 3640
rect 1100 3580 1300 3600
use diff_pair  diff_pair_0
timestamp 1730311536
transform 1 0 -234 0 1 2300
box 234 -2300 2665 1550
use sky130_fd_pr__pfet_01v8_J24L55  sky130_fd_pr__pfet_01v8_J24L55_0
timestamp 1730316371
transform 0 1 1200 -1 0 4794
box -194 -200 194 200
<< end >>
