magic
tech sky130A
magscale 1 2
timestamp 1731631080
<< xpolycontact >>
rect 297 4104 367 4536
rect -367 -4536 -297 -4104
<< xpolyres >>
rect -367 3930 -131 4000
rect -367 -4104 -297 3930
rect -201 -3930 -131 3930
rect -35 3930 201 4000
rect -35 -3930 35 3930
rect -201 -4000 35 -3930
rect 131 -3930 201 3930
rect 297 -3930 367 4104
rect 131 -4000 367 -3930
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 40 m 1 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 1.151meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_0p35_UYKEAK parameters
<< end >>
