magic
tech sky130A
magscale 1 2
timestamp 1730605901
<< xpolycontact >>
rect -573 7984 573 8416
rect -573 -8416 573 -7984
<< xpolyres >>
rect -573 -7984 573 7984
<< viali >>
rect -557 8001 557 8398
rect -557 -8398 557 -8001
<< metal1 >>
rect -569 8398 569 8404
rect -569 8001 -557 8398
rect 557 8001 569 8398
rect -569 7995 569 8001
rect -569 -8001 569 -7995
rect -569 -8398 -557 -8001
rect 557 -8398 569 -8001
rect -569 -8404 569 -8398
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 80.0 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 27.988k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_5p73_6QC7Y6 parameters
<< end >>
