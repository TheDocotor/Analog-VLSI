magic
tech sky130A
magscale 1 2
timestamp 1731632322
<< nmos >>
rect -100 -969 100 1031
<< ndiff >>
rect -158 1019 -100 1031
rect -158 -957 -146 1019
rect -112 -957 -100 1019
rect -158 -969 -100 -957
rect 100 1019 158 1031
rect 100 -957 112 1019
rect 146 -957 158 1019
rect 100 -969 158 -957
<< ndiffc >>
rect -146 -957 -112 1019
rect 112 -957 146 1019
<< poly >>
rect -100 1031 100 1057
rect -100 -1007 100 -969
rect -100 -1041 -84 -1007
rect 84 -1041 100 -1007
rect -100 -1057 100 -1041
<< polycont >>
rect -84 -1041 84 -1007
<< locali >>
rect -146 1019 -112 1035
rect -146 -973 -112 -957
rect 112 1019 146 1035
rect 112 -973 146 -957
rect -100 -1041 -84 -1007
rect 84 -1041 100 -1007
<< viali >>
rect -146 -957 -112 1019
rect 112 -957 146 1019
rect -84 -1041 84 -1007
<< metal1 >>
rect -152 1019 -106 1031
rect -152 -957 -146 1019
rect -112 -957 -106 1019
rect -152 -969 -106 -957
rect 106 1019 152 1031
rect 106 -957 112 1019
rect 146 -957 152 1019
rect 106 -969 152 -957
rect -96 -1007 96 -1001
rect -96 -1041 -84 -1007
rect 84 -1041 96 -1007
rect -96 -1047 96 -1041
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_7JY9FK parameters
<< end >>
