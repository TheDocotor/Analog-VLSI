magic
tech sky130A
magscale 1 2
timestamp 1732735281
<< nwell >>
rect -4480 -760 -680 40
<< pmos >>
rect -4100 -120 -900 -80
rect -4100 -240 -900 -200
rect -4100 -360 -900 -320
rect -4100 -480 -900 -440
rect -4100 -600 -900 -560
<< pdiff >>
rect -4100 -20 -900 0
rect -4100 -60 -4080 -20
rect -920 -60 -900 -20
rect -4100 -80 -900 -60
rect -4100 -140 -900 -120
rect -4100 -180 -4080 -140
rect -920 -180 -900 -140
rect -4100 -200 -900 -180
rect -4100 -260 -900 -240
rect -4100 -300 -4080 -260
rect -920 -300 -900 -260
rect -4100 -320 -900 -300
rect -4100 -380 -900 -360
rect -4100 -420 -4080 -380
rect -920 -420 -900 -380
rect -4100 -440 -900 -420
rect -4100 -500 -900 -480
rect -4100 -540 -4080 -500
rect -920 -540 -900 -500
rect -4100 -560 -900 -540
rect -4100 -620 -900 -600
rect -4100 -660 -4080 -620
rect -920 -660 -900 -620
rect -4100 -680 -900 -660
<< pdiffc >>
rect -4080 -60 -920 -20
rect -4080 -180 -920 -140
rect -4080 -300 -920 -260
rect -4080 -420 -920 -380
rect -4080 -540 -920 -500
rect -4080 -660 -920 -620
<< poly >>
rect -4440 -120 -4100 -80
rect -900 -120 -800 -80
rect -4440 -560 -4400 -120
rect -4320 -200 -4280 -120
rect -4320 -240 -4100 -200
rect -900 -240 -800 -200
rect -4320 -320 -4280 -240
rect -4320 -360 -4100 -320
rect -900 -360 -800 -320
rect -4320 -440 -4280 -360
rect -4320 -480 -4100 -440
rect -900 -480 -800 -440
rect -4320 -560 -4280 -480
rect -4440 -600 -4100 -560
rect -900 -600 -800 -560
<< polycont >>
rect -4400 -560 -4320 -120
<< locali >>
rect -4240 -20 -900 0
rect -4240 -60 -4080 -20
rect -920 -60 -900 -20
rect -4240 -80 -900 -60
rect -4440 -120 -4280 -80
rect -4440 -560 -4400 -120
rect -4320 -560 -4280 -120
rect -4240 -240 -4200 -80
rect -4100 -140 -720 -120
rect -4100 -180 -4080 -140
rect -920 -180 -720 -140
rect -4100 -200 -720 -180
rect -4240 -260 -900 -240
rect -4240 -300 -4080 -260
rect -920 -300 -900 -260
rect -4240 -320 -900 -300
rect -4240 -480 -4200 -320
rect -800 -360 -720 -200
rect -4100 -380 -720 -360
rect -4100 -420 -4080 -380
rect -920 -420 -720 -380
rect -4100 -440 -720 -420
rect -4240 -500 -900 -480
rect -4240 -540 -4080 -500
rect -920 -540 -900 -500
rect -4240 -560 -900 -540
rect -4440 -600 -4280 -560
rect -800 -600 -720 -440
rect -4100 -620 -720 -600
rect -4100 -660 -4080 -620
rect -920 -660 -720 -620
rect -4100 -680 -720 -660
<< labels >>
flabel pdiffc -2479 -44 -2479 -44 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont -4361 -336 -4361 -336 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel pdiffc -2475 -645 -2475 -645 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell -4367 -19 -4367 -19 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
