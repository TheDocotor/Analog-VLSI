magic
tech sky130A
magscale 1 2
timestamp 1729559727
use sky130_fd_pr__res_xhigh_po_0p69_C432MY  sky130_fd_pr__res_xhigh_po_0p69_C432MY_0
timestamp 1729559727
transform 1 0 16 0 1 674
box -69 -727 69 727
<< end >>
