magic
tech sky130A
magscale 1 2
timestamp 1730605901
<< nwell >>
rect 2475 450 3975 1650
<< pmos >>
rect 2900 1400 3700 1500
rect 2900 1200 3700 1300
rect 2900 1000 3700 1100
rect 2900 800 3700 900
rect 2900 600 3700 700
<< pdiff >>
rect 2900 1575 3700 1600
rect 2900 1525 2925 1575
rect 3675 1525 3700 1575
rect 2900 1500 3700 1525
rect 2900 1375 3700 1400
rect 2900 1325 2925 1375
rect 3675 1325 3700 1375
rect 2900 1300 3700 1325
rect 2900 1175 3700 1200
rect 2900 1125 2925 1175
rect 3675 1125 3700 1175
rect 2900 1100 3700 1125
rect 2900 975 3700 1000
rect 2900 925 2925 975
rect 3675 925 3700 975
rect 2900 900 3700 925
rect 2900 775 3700 800
rect 2900 725 2925 775
rect 3675 725 3700 775
rect 2900 700 3700 725
rect 2900 575 3700 600
rect 2900 525 2925 575
rect 3675 525 3700 575
rect 2900 500 3700 525
<< pdiffc >>
rect 2925 1525 3675 1575
rect 2925 1325 3675 1375
rect 2925 1125 3675 1175
rect 2925 925 3675 975
rect 2925 725 3675 775
rect 2925 525 3675 575
<< poly >>
rect 2500 1475 2900 1500
rect 2500 625 2525 1475
rect 2575 1400 2900 1475
rect 3700 1400 3900 1500
rect 2575 1300 2650 1400
rect 2575 1200 2900 1300
rect 3700 1200 3900 1300
rect 2575 1100 2650 1200
rect 2575 1000 2900 1100
rect 3700 1000 3900 1100
rect 2575 900 2650 1000
rect 2575 800 2900 900
rect 3700 800 3900 900
rect 2575 700 2650 800
rect 2575 625 2900 700
rect 2500 600 2900 625
rect 3700 600 3900 700
<< polycont >>
rect 2525 625 2575 1475
<< locali >>
rect 2650 1575 3800 1600
rect 2650 1525 2925 1575
rect 3675 1525 3800 1575
rect 2650 1500 3800 1525
rect 2500 1475 2600 1500
rect 2500 625 2525 1475
rect 2575 625 2600 1475
rect 2650 1200 2750 1500
rect 3850 1400 3950 1500
rect 2800 1375 3950 1400
rect 2800 1325 2925 1375
rect 3675 1325 3950 1375
rect 2800 1300 3950 1325
rect 2650 1175 3800 1200
rect 2650 1125 2925 1175
rect 3675 1125 3800 1175
rect 2650 1100 3800 1125
rect 2650 800 2750 1100
rect 3850 1000 3950 1300
rect 2800 975 3950 1000
rect 2800 925 2925 975
rect 3675 925 3950 975
rect 2800 900 3950 925
rect 2650 775 3800 800
rect 2650 725 2925 775
rect 3675 725 3800 775
rect 2650 700 3800 725
rect 2500 600 2600 625
rect 3850 600 3950 900
rect 2800 575 3950 600
rect 2800 525 2925 575
rect 3675 525 3950 575
rect 2800 500 3950 525
<< labels >>
flabel pdiffc 3300 1550 3300 1550 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont 2550 1050 2550 1050 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel pdiffc 3325 550 3325 550 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell 2550 1575 2550 1575 0 FreeSans 800 0 0 0 B
port 3 nsew
<< properties >>
string p20x05 parameters
<< end >>
