magic
tech sky130A
magscale 1 2
timestamp 1730302828
<< nwell >>
rect -25 -1150 1075 550
<< pmos >>
rect 300 200 900 400
rect 300 -100 900 100
rect 300 -400 900 -200
rect 300 -700 900 -500
rect 300 -1000 900 -800
<< pdiff >>
rect 300 475 900 500
rect 300 425 325 475
rect 875 425 900 475
rect 300 400 900 425
rect 300 175 900 200
rect 300 125 325 175
rect 875 125 900 175
rect 300 100 900 125
rect 300 -125 900 -100
rect 300 -175 325 -125
rect 875 -175 900 -125
rect 300 -200 900 -175
rect 300 -425 900 -400
rect 300 -475 325 -425
rect 875 -475 900 -425
rect 300 -500 900 -475
rect 300 -725 900 -700
rect 300 -775 325 -725
rect 875 -775 900 -725
rect 300 -800 900 -775
rect 300 -1025 900 -1000
rect 300 -1075 325 -1025
rect 875 -1075 900 -1025
rect 300 -1100 900 -1075
<< pdiffc >>
rect 325 425 875 475
rect 325 125 875 175
rect 325 -175 875 -125
rect 325 -475 875 -425
rect 325 -775 875 -725
rect 325 -1075 875 -1025
<< poly >>
rect 0 375 200 400
rect 0 -975 25 375
rect 75 100 200 375
rect 250 200 300 400
rect 900 200 1000 400
rect 75 -100 300 100
rect 900 -100 1000 100
rect 75 -200 200 -100
rect 75 -400 300 -200
rect 900 -400 1000 -200
rect 75 -500 200 -400
rect 75 -700 300 -500
rect 900 -700 1000 -500
rect 75 -800 200 -700
rect 75 -975 300 -800
rect 0 -1000 300 -975
rect 900 -1000 1000 -800
<< polycont >>
rect 25 -975 75 375
<< locali >>
rect 150 475 900 500
rect 150 425 325 475
rect 875 425 900 475
rect 150 400 900 425
rect 0 375 100 400
rect 0 -975 25 375
rect 75 -975 100 375
rect 150 -100 250 400
rect 300 175 1050 200
rect 300 125 325 175
rect 875 125 1050 175
rect 300 100 1050 125
rect 150 -125 900 -100
rect 150 -175 325 -125
rect 875 -175 900 -125
rect 150 -200 900 -175
rect 150 -700 250 -200
rect 950 -400 1050 100
rect 300 -425 1050 -400
rect 300 -475 325 -425
rect 875 -475 1050 -425
rect 300 -500 1050 -475
rect 150 -725 900 -700
rect 150 -775 325 -725
rect 875 -775 900 -725
rect 150 -800 900 -775
rect 0 -1000 100 -975
rect 950 -1000 1050 -500
rect 300 -1025 1050 -1000
rect 300 -1075 325 -1025
rect 875 -1075 1050 -1025
rect 300 -1100 1050 -1075
<< labels >>
flabel pdiffc 600 450 600 450 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont 50 -300 50 -300 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel pdiffc 625 -1050 625 -1050 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell 50 475 50 475 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
