magic
tech sky130A
magscale 1 2
timestamp 1729093895
<< pwell >>
rect -1400 200 0 2600
<< nmos >>
rect -1220 400 -1000 2400
rect -940 400 -720 2400
rect -660 400 -440 2400
rect -380 400 -160 2400
<< ndiff >>
rect -1280 2380 -1220 2400
rect -1280 420 -1265 2380
rect -1231 420 -1220 2380
rect -1280 400 -1220 420
rect -1000 2380 -940 2400
rect -1000 420 -985 2380
rect -951 420 -940 2380
rect -1000 400 -940 420
rect -720 2380 -660 2400
rect -720 420 -705 2380
rect -671 420 -660 2380
rect -720 400 -660 420
rect -440 2380 -380 2400
rect -440 420 -425 2380
rect -391 420 -380 2380
rect -440 400 -380 420
rect -160 2380 -100 2400
rect -160 420 -145 2380
rect -111 420 -100 2380
rect -160 400 -100 420
<< ndiffc >>
rect -1265 420 -1231 2380
rect -985 420 -951 2380
rect -705 420 -671 2380
rect -425 420 -391 2380
rect -145 420 -111 2380
<< poly >>
rect -1220 2560 -160 2580
rect -1220 2520 -1180 2560
rect -200 2520 -160 2560
rect -1220 2500 -160 2520
rect -1220 2400 -1000 2500
rect -940 2400 -720 2500
rect -660 2400 -440 2500
rect -380 2400 -160 2500
rect -1220 300 -1000 400
rect -940 300 -720 400
rect -660 300 -440 400
rect -380 300 -160 400
<< polycont >>
rect -1180 2520 -200 2560
<< locali >>
rect -1220 2520 -1180 2560
rect -200 2520 -160 2560
rect -1270 2440 -110 2480
rect -1270 2380 -1230 2440
rect -1270 420 -1265 2380
rect -1231 420 -1230 2380
rect -1270 395 -1230 420
rect -990 2380 -950 2405
rect -990 420 -985 2380
rect -951 420 -950 2380
rect -990 290 -950 420
rect -710 2380 -670 2440
rect -710 420 -705 2380
rect -671 420 -670 2380
rect -710 395 -670 420
rect -430 2380 -390 2405
rect -430 420 -425 2380
rect -391 420 -390 2380
rect -430 290 -390 420
rect -150 2380 -110 2440
rect -150 420 -145 2380
rect -111 420 -110 2380
rect -150 395 -110 420
rect -990 250 -390 290
<< viali >>
rect -1180 2520 -200 2560
rect -1265 420 -1231 2380
rect -985 420 -951 2380
rect -705 420 -671 2380
rect -425 420 -391 2380
rect -145 420 -111 2380
<< metal1 >>
rect -1190 2560 -190 2570
rect -1220 2520 -1180 2560
rect -200 2520 -160 2560
rect -1190 2510 -190 2520
rect -1275 2380 -1225 2400
rect -1275 420 -1265 2380
rect -1231 420 -1225 2380
rect -1275 400 -1225 420
rect -995 2380 -945 2400
rect -995 420 -985 2380
rect -951 420 -945 2380
rect -995 400 -945 420
rect -715 2380 -665 2400
rect -715 420 -705 2380
rect -671 420 -665 2380
rect -715 400 -665 420
rect -435 2380 -385 2400
rect -435 420 -425 2380
rect -391 420 -385 2380
rect -435 400 -385 420
rect -155 2380 -105 2400
rect -155 420 -145 2380
rect -111 420 -105 2380
rect -155 400 -105 420
<< labels >>
flabel viali -744 2540 -744 2540 0 FreeSans 800 0 0 0 G
port 2 nsew
flabel locali -141 2450 -141 2450 0 FreeSans 800 0 0 0 S
port 3 nsew
flabel locali -683 266 -683 266 0 FreeSans 800 0 0 0 D
port 1 nsew
flabel pwell -39 1659 -39 1659 0 FreeSans 800 0 0 0 B
port 4 nsew
<< end >>
