* SPICE3 file created from pmos.ext - technology: sky130A

X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.27 pd=2.4 as=0.27 ps=2.4 w=0.9 l=1
