** sch_path: /home/renslow/Documents/ece5120/hw03/mag/nmos_tb.sch
**.subckt nmos_tb
Vd1 D1v8 D 0
.save i(vd1)
x1 D G1v8 S B nmos_40
**** begin user architecture code

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
.include /home/renslow/Documents/ece5120/hw03/mag/nmos_40.spice
vg G1v8 0 1.8
vs s 0 0
vd D1v8 0 1.8
vb b 0 0
.control
save all

dc vd 0 1.8 0.005 vg 0 1.8 0.1
write my_nmos_tb.raw

plot all.vd1#branch vs D1v8
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/magic/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/magic/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/magic/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/magic/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.end
