magic
tech sky130A
magscale 1 2
timestamp 1732734633
<< nwell >>
rect -10800 -9960 6000 -120
<< pmos >>
rect -10300 -320 5700 -280
rect -10300 -440 5700 -400
rect -10300 -560 5700 -520
rect -10300 -680 5700 -640
rect -10300 -800 5700 -760
rect -10300 -920 5700 -880
rect -10300 -1040 5700 -1000
rect -10300 -1160 5700 -1120
rect -10300 -1280 5700 -1240
rect -10300 -1400 5700 -1360
rect -10300 -1520 5700 -1480
rect -10300 -1640 5700 -1600
rect -10300 -1760 5700 -1720
rect -10300 -1880 5700 -1840
rect -10300 -2000 5700 -1960
rect -10300 -2120 5700 -2080
rect -10300 -2240 5700 -2200
rect -10300 -2360 5700 -2320
rect -10300 -2480 5700 -2440
rect -10300 -2600 5700 -2560
rect -10300 -2720 5700 -2680
rect -10300 -2840 5700 -2800
rect -10300 -2960 5700 -2920
rect -10300 -3080 5700 -3040
rect -10300 -3200 5700 -3160
rect -10300 -3320 5700 -3280
rect -10300 -3440 5700 -3400
rect -10300 -3560 5700 -3520
rect -10300 -3680 5700 -3640
rect -10300 -3800 5700 -3760
rect -10300 -3920 5700 -3880
rect -10300 -4040 5700 -4000
rect -10300 -4160 5700 -4120
rect -10300 -4280 5700 -4240
rect -10300 -4400 5700 -4360
rect -10300 -4520 5700 -4480
rect -10300 -4640 5700 -4600
rect -10300 -4760 5700 -4720
rect -10300 -4880 5700 -4840
rect -10300 -5000 5700 -4960
rect -10300 -5120 5700 -5080
rect -10300 -5240 5700 -5200
rect -10300 -5360 5700 -5320
rect -10300 -5480 5700 -5440
rect -10300 -5600 5700 -5560
rect -10300 -5720 5700 -5680
rect -10300 -5840 5700 -5800
rect -10300 -5960 5700 -5920
rect -10300 -6080 5700 -6040
rect -10300 -6200 5700 -6160
rect -10300 -6320 5700 -6280
rect -10300 -6440 5700 -6400
rect -10300 -6560 5700 -6520
rect -10300 -6680 5700 -6640
rect -10300 -6800 5700 -6760
rect -10300 -6920 5700 -6880
rect -10300 -7040 5700 -7000
rect -10300 -7160 5700 -7120
rect -10300 -7280 5700 -7240
rect -10300 -7400 5700 -7360
rect -10300 -7520 5700 -7480
rect -10300 -7640 5700 -7600
rect -10300 -7760 5700 -7720
rect -10300 -7880 5700 -7840
rect -10300 -8000 5700 -7960
rect -10300 -8120 5700 -8080
rect -10300 -8240 5700 -8200
rect -10300 -8360 5700 -8320
rect -10300 -8480 5700 -8440
rect -10300 -8600 5700 -8560
rect -10300 -8720 5700 -8680
rect -10300 -8840 5700 -8800
rect -10300 -8960 5700 -8920
rect -10300 -9080 5700 -9040
rect -10300 -9200 5700 -9160
rect -10300 -9320 5700 -9280
rect -10300 -9440 5700 -9400
rect -10300 -9560 5700 -9520
rect -10300 -9680 5700 -9640
rect -10300 -9800 5700 -9760
<< pdiff >>
rect -10300 -220 5700 -200
rect -10300 -260 -10280 -220
rect 5680 -260 5700 -220
rect -10300 -280 5700 -260
rect -10300 -340 5700 -320
rect -10300 -380 -10280 -340
rect 5680 -380 5700 -340
rect -10300 -400 5700 -380
rect -10300 -460 5700 -440
rect -10300 -500 -10280 -460
rect 5680 -500 5700 -460
rect -10300 -520 5700 -500
rect -10300 -580 5700 -560
rect -10300 -620 -10280 -580
rect 5680 -620 5700 -580
rect -10300 -640 5700 -620
rect -10300 -700 5700 -680
rect -10300 -740 -10280 -700
rect 5680 -740 5700 -700
rect -10300 -760 5700 -740
rect -10300 -820 5700 -800
rect -10300 -860 -10280 -820
rect 5680 -860 5700 -820
rect -10300 -880 5700 -860
rect -10300 -940 5700 -920
rect -10300 -980 -10280 -940
rect 5680 -980 5700 -940
rect -10300 -1000 5700 -980
rect -10300 -1060 5700 -1040
rect -10300 -1100 -10280 -1060
rect 5680 -1100 5700 -1060
rect -10300 -1120 5700 -1100
rect -10300 -1180 5700 -1160
rect -10300 -1220 -10280 -1180
rect 5680 -1220 5700 -1180
rect -10300 -1240 5700 -1220
rect -10300 -1300 5700 -1280
rect -10300 -1340 -10280 -1300
rect 5680 -1340 5700 -1300
rect -10300 -1360 5700 -1340
rect -10300 -1420 5700 -1400
rect -10300 -1460 -10280 -1420
rect 5680 -1460 5700 -1420
rect -10300 -1480 5700 -1460
rect -10300 -1540 5700 -1520
rect -10300 -1580 -10280 -1540
rect 5680 -1580 5700 -1540
rect -10300 -1600 5700 -1580
rect -10300 -1660 5700 -1640
rect -10300 -1700 -10280 -1660
rect 5680 -1700 5700 -1660
rect -10300 -1720 5700 -1700
rect -10300 -1780 5700 -1760
rect -10300 -1820 -10280 -1780
rect 5680 -1820 5700 -1780
rect -10300 -1840 5700 -1820
rect -10300 -1900 5700 -1880
rect -10300 -1940 -10280 -1900
rect 5680 -1940 5700 -1900
rect -10300 -1960 5700 -1940
rect -10300 -2020 5700 -2000
rect -10300 -2060 -10280 -2020
rect 5680 -2060 5700 -2020
rect -10300 -2080 5700 -2060
rect -10300 -2140 5700 -2120
rect -10300 -2180 -10280 -2140
rect 5680 -2180 5700 -2140
rect -10300 -2200 5700 -2180
rect -10300 -2260 5700 -2240
rect -10300 -2300 -10280 -2260
rect 5680 -2300 5700 -2260
rect -10300 -2320 5700 -2300
rect -10300 -2380 5700 -2360
rect -10300 -2420 -10280 -2380
rect 5680 -2420 5700 -2380
rect -10300 -2440 5700 -2420
rect -10300 -2500 5700 -2480
rect -10300 -2540 -10280 -2500
rect 5680 -2540 5700 -2500
rect -10300 -2560 5700 -2540
rect -10300 -2620 5700 -2600
rect -10300 -2660 -10280 -2620
rect 5680 -2660 5700 -2620
rect -10300 -2680 5700 -2660
rect -10300 -2740 5700 -2720
rect -10300 -2780 -10280 -2740
rect 5680 -2780 5700 -2740
rect -10300 -2800 5700 -2780
rect -10300 -2860 5700 -2840
rect -10300 -2900 -10280 -2860
rect 5680 -2900 5700 -2860
rect -10300 -2920 5700 -2900
rect -10300 -2980 5700 -2960
rect -10300 -3020 -10280 -2980
rect 5680 -3020 5700 -2980
rect -10300 -3040 5700 -3020
rect -10300 -3100 5700 -3080
rect -10300 -3140 -10280 -3100
rect 5680 -3140 5700 -3100
rect -10300 -3160 5700 -3140
rect -10300 -3220 5700 -3200
rect -10300 -3260 -10280 -3220
rect 5680 -3260 5700 -3220
rect -10300 -3280 5700 -3260
rect -10300 -3340 5700 -3320
rect -10300 -3380 -10280 -3340
rect 5680 -3380 5700 -3340
rect -10300 -3400 5700 -3380
rect -10300 -3460 5700 -3440
rect -10300 -3500 -10280 -3460
rect 5680 -3500 5700 -3460
rect -10300 -3520 5700 -3500
rect -10300 -3580 5700 -3560
rect -10300 -3620 -10280 -3580
rect 5680 -3620 5700 -3580
rect -10300 -3640 5700 -3620
rect -10300 -3700 5700 -3680
rect -10300 -3740 -10280 -3700
rect 5680 -3740 5700 -3700
rect -10300 -3760 5700 -3740
rect -10300 -3820 5700 -3800
rect -10300 -3860 -10280 -3820
rect 5680 -3860 5700 -3820
rect -10300 -3880 5700 -3860
rect -10300 -3940 5700 -3920
rect -10300 -3980 -10280 -3940
rect 5680 -3980 5700 -3940
rect -10300 -4000 5700 -3980
rect -10300 -4060 5700 -4040
rect -10300 -4100 -10280 -4060
rect 5680 -4100 5700 -4060
rect -10300 -4120 5700 -4100
rect -10300 -4180 5700 -4160
rect -10300 -4220 -10280 -4180
rect 5680 -4220 5700 -4180
rect -10300 -4240 5700 -4220
rect -10300 -4300 5700 -4280
rect -10300 -4340 -10280 -4300
rect 5680 -4340 5700 -4300
rect -10300 -4360 5700 -4340
rect -10300 -4420 5700 -4400
rect -10300 -4460 -10280 -4420
rect 5680 -4460 5700 -4420
rect -10300 -4480 5700 -4460
rect -10300 -4540 5700 -4520
rect -10300 -4580 -10280 -4540
rect 5680 -4580 5700 -4540
rect -10300 -4600 5700 -4580
rect -10300 -4660 5700 -4640
rect -10300 -4700 -10280 -4660
rect 5680 -4700 5700 -4660
rect -10300 -4720 5700 -4700
rect -10300 -4780 5700 -4760
rect -10300 -4820 -10280 -4780
rect 5680 -4820 5700 -4780
rect -10300 -4840 5700 -4820
rect -10300 -4900 5700 -4880
rect -10300 -4940 -10280 -4900
rect 5680 -4940 5700 -4900
rect -10300 -4960 5700 -4940
rect -10300 -5020 5700 -5000
rect -10300 -5060 -10280 -5020
rect 5680 -5060 5700 -5020
rect -10300 -5080 5700 -5060
rect -10300 -5140 5700 -5120
rect -10300 -5180 -10280 -5140
rect 5680 -5180 5700 -5140
rect -10300 -5200 5700 -5180
rect -10300 -5260 5700 -5240
rect -10300 -5300 -10280 -5260
rect 5680 -5300 5700 -5260
rect -10300 -5320 5700 -5300
rect -10300 -5380 5700 -5360
rect -10300 -5420 -10280 -5380
rect 5680 -5420 5700 -5380
rect -10300 -5440 5700 -5420
rect -10300 -5500 5700 -5480
rect -10300 -5540 -10280 -5500
rect 5680 -5540 5700 -5500
rect -10300 -5560 5700 -5540
rect -10300 -5620 5700 -5600
rect -10300 -5660 -10280 -5620
rect 5680 -5660 5700 -5620
rect -10300 -5680 5700 -5660
rect -10300 -5740 5700 -5720
rect -10300 -5780 -10280 -5740
rect 5680 -5780 5700 -5740
rect -10300 -5800 5700 -5780
rect -10300 -5860 5700 -5840
rect -10300 -5900 -10280 -5860
rect 5680 -5900 5700 -5860
rect -10300 -5920 5700 -5900
rect -10300 -5980 5700 -5960
rect -10300 -6020 -10280 -5980
rect 5680 -6020 5700 -5980
rect -10300 -6040 5700 -6020
rect -10300 -6100 5700 -6080
rect -10300 -6140 -10280 -6100
rect 5680 -6140 5700 -6100
rect -10300 -6160 5700 -6140
rect -10300 -6220 5700 -6200
rect -10300 -6260 -10280 -6220
rect 5680 -6260 5700 -6220
rect -10300 -6280 5700 -6260
rect -10300 -6340 5700 -6320
rect -10300 -6380 -10280 -6340
rect 5680 -6380 5700 -6340
rect -10300 -6400 5700 -6380
rect -10300 -6460 5700 -6440
rect -10300 -6500 -10280 -6460
rect 5680 -6500 5700 -6460
rect -10300 -6520 5700 -6500
rect -10300 -6580 5700 -6560
rect -10300 -6620 -10280 -6580
rect 5680 -6620 5700 -6580
rect -10300 -6640 5700 -6620
rect -10300 -6700 5700 -6680
rect -10300 -6740 -10280 -6700
rect 5680 -6740 5700 -6700
rect -10300 -6760 5700 -6740
rect -10300 -6820 5700 -6800
rect -10300 -6860 -10280 -6820
rect 5680 -6860 5700 -6820
rect -10300 -6880 5700 -6860
rect -10300 -6940 5700 -6920
rect -10300 -6980 -10280 -6940
rect 5680 -6980 5700 -6940
rect -10300 -7000 5700 -6980
rect -10300 -7060 5700 -7040
rect -10300 -7100 -10280 -7060
rect 5680 -7100 5700 -7060
rect -10300 -7120 5700 -7100
rect -10300 -7180 5700 -7160
rect -10300 -7220 -10280 -7180
rect 5680 -7220 5700 -7180
rect -10300 -7240 5700 -7220
rect -10300 -7300 5700 -7280
rect -10300 -7340 -10280 -7300
rect 5680 -7340 5700 -7300
rect -10300 -7360 5700 -7340
rect -10300 -7420 5700 -7400
rect -10300 -7460 -10280 -7420
rect 5680 -7460 5700 -7420
rect -10300 -7480 5700 -7460
rect -10300 -7540 5700 -7520
rect -10300 -7580 -10280 -7540
rect 5680 -7580 5700 -7540
rect -10300 -7600 5700 -7580
rect -10300 -7660 5700 -7640
rect -10300 -7700 -10280 -7660
rect 5680 -7700 5700 -7660
rect -10300 -7720 5700 -7700
rect -10300 -7780 5700 -7760
rect -10300 -7820 -10280 -7780
rect 5680 -7820 5700 -7780
rect -10300 -7840 5700 -7820
rect -10300 -7900 5700 -7880
rect -10300 -7940 -10280 -7900
rect 5680 -7940 5700 -7900
rect -10300 -7960 5700 -7940
rect -10300 -8020 5700 -8000
rect -10300 -8060 -10280 -8020
rect 5680 -8060 5700 -8020
rect -10300 -8080 5700 -8060
rect -10300 -8140 5700 -8120
rect -10300 -8180 -10280 -8140
rect 5680 -8180 5700 -8140
rect -10300 -8200 5700 -8180
rect -10300 -8260 5700 -8240
rect -10300 -8300 -10280 -8260
rect 5680 -8300 5700 -8260
rect -10300 -8320 5700 -8300
rect -10300 -8380 5700 -8360
rect -10300 -8420 -10280 -8380
rect 5680 -8420 5700 -8380
rect -10300 -8440 5700 -8420
rect -10300 -8500 5700 -8480
rect -10300 -8540 -10280 -8500
rect 5680 -8540 5700 -8500
rect -10300 -8560 5700 -8540
rect -10300 -8620 5700 -8600
rect -10300 -8660 -10280 -8620
rect 5680 -8660 5700 -8620
rect -10300 -8680 5700 -8660
rect -10300 -8740 5700 -8720
rect -10300 -8780 -10280 -8740
rect 5680 -8780 5700 -8740
rect -10300 -8800 5700 -8780
rect -10300 -8860 5700 -8840
rect -10300 -8900 -10280 -8860
rect 5680 -8900 5700 -8860
rect -10300 -8920 5700 -8900
rect -10300 -8980 5700 -8960
rect -10300 -9020 -10280 -8980
rect 5680 -9020 5700 -8980
rect -10300 -9040 5700 -9020
rect -10300 -9100 5700 -9080
rect -10300 -9140 -10280 -9100
rect 5680 -9140 5700 -9100
rect -10300 -9160 5700 -9140
rect -10300 -9220 5700 -9200
rect -10300 -9260 -10280 -9220
rect 5680 -9260 5700 -9220
rect -10300 -9280 5700 -9260
rect -10300 -9340 5700 -9320
rect -10300 -9380 -10280 -9340
rect 5680 -9380 5700 -9340
rect -10300 -9400 5700 -9380
rect -10300 -9460 5700 -9440
rect -10300 -9500 -10280 -9460
rect 5680 -9500 5700 -9460
rect -10300 -9520 5700 -9500
rect -10300 -9580 5700 -9560
rect -10300 -9620 -10280 -9580
rect 5680 -9620 5700 -9580
rect -10300 -9640 5700 -9620
rect -10300 -9700 5700 -9680
rect -10300 -9740 -10280 -9700
rect 5680 -9740 5700 -9700
rect -10300 -9760 5700 -9740
rect -10300 -9820 5700 -9800
rect -10300 -9860 -10280 -9820
rect 5680 -9860 5700 -9820
rect -10300 -9880 5700 -9860
<< pdiffc >>
rect -10280 -260 5680 -220
rect -10280 -380 5680 -340
rect -10280 -500 5680 -460
rect -10280 -620 5680 -580
rect -10280 -740 5680 -700
rect -10280 -860 5680 -820
rect -10280 -980 5680 -940
rect -10280 -1100 5680 -1060
rect -10280 -1220 5680 -1180
rect -10280 -1340 5680 -1300
rect -10280 -1460 5680 -1420
rect -10280 -1580 5680 -1540
rect -10280 -1700 5680 -1660
rect -10280 -1820 5680 -1780
rect -10280 -1940 5680 -1900
rect -10280 -2060 5680 -2020
rect -10280 -2180 5680 -2140
rect -10280 -2300 5680 -2260
rect -10280 -2420 5680 -2380
rect -10280 -2540 5680 -2500
rect -10280 -2660 5680 -2620
rect -10280 -2780 5680 -2740
rect -10280 -2900 5680 -2860
rect -10280 -3020 5680 -2980
rect -10280 -3140 5680 -3100
rect -10280 -3260 5680 -3220
rect -10280 -3380 5680 -3340
rect -10280 -3500 5680 -3460
rect -10280 -3620 5680 -3580
rect -10280 -3740 5680 -3700
rect -10280 -3860 5680 -3820
rect -10280 -3980 5680 -3940
rect -10280 -4100 5680 -4060
rect -10280 -4220 5680 -4180
rect -10280 -4340 5680 -4300
rect -10280 -4460 5680 -4420
rect -10280 -4580 5680 -4540
rect -10280 -4700 5680 -4660
rect -10280 -4820 5680 -4780
rect -10280 -4940 5680 -4900
rect -10280 -5060 5680 -5020
rect -10280 -5180 5680 -5140
rect -10280 -5300 5680 -5260
rect -10280 -5420 5680 -5380
rect -10280 -5540 5680 -5500
rect -10280 -5660 5680 -5620
rect -10280 -5780 5680 -5740
rect -10280 -5900 5680 -5860
rect -10280 -6020 5680 -5980
rect -10280 -6140 5680 -6100
rect -10280 -6260 5680 -6220
rect -10280 -6380 5680 -6340
rect -10280 -6500 5680 -6460
rect -10280 -6620 5680 -6580
rect -10280 -6740 5680 -6700
rect -10280 -6860 5680 -6820
rect -10280 -6980 5680 -6940
rect -10280 -7100 5680 -7060
rect -10280 -7220 5680 -7180
rect -10280 -7340 5680 -7300
rect -10280 -7460 5680 -7420
rect -10280 -7580 5680 -7540
rect -10280 -7700 5680 -7660
rect -10280 -7820 5680 -7780
rect -10280 -7940 5680 -7900
rect -10280 -8060 5680 -8020
rect -10280 -8180 5680 -8140
rect -10280 -8300 5680 -8260
rect -10280 -8420 5680 -8380
rect -10280 -8540 5680 -8500
rect -10280 -8660 5680 -8620
rect -10280 -8780 5680 -8740
rect -10280 -8900 5680 -8860
rect -10280 -9020 5680 -8980
rect -10280 -9140 5680 -9100
rect -10280 -9260 5680 -9220
rect -10280 -9380 5680 -9340
rect -10280 -9500 5680 -9460
rect -10280 -9620 5680 -9580
rect -10280 -9740 5680 -9700
rect -10280 -9860 5680 -9820
<< poly >>
rect -10680 -320 -10300 -280
rect 5700 -320 5800 -280
rect -10680 -9760 -10640 -320
rect -10600 -400 -10560 -320
rect -10600 -440 -10300 -400
rect 5700 -440 5800 -400
rect -10600 -520 -10560 -440
rect -10600 -560 -10300 -520
rect 5700 -560 5800 -520
rect -10600 -640 -10560 -560
rect -10600 -680 -10300 -640
rect 5700 -680 5800 -640
rect -10600 -760 -10560 -680
rect -10600 -800 -10300 -760
rect 5700 -800 5800 -760
rect -10600 -880 -10560 -800
rect -10600 -920 -10300 -880
rect 5700 -920 5800 -880
rect -10600 -1000 -10560 -920
rect -10600 -1040 -10300 -1000
rect 5700 -1040 5800 -1000
rect -10600 -1120 -10560 -1040
rect -10600 -1160 -10300 -1120
rect 5700 -1160 5800 -1120
rect -10600 -1240 -10560 -1160
rect -10600 -1280 -10300 -1240
rect 5700 -1280 5800 -1240
rect -10600 -1360 -10560 -1280
rect -10600 -1400 -10300 -1360
rect 5700 -1400 5800 -1360
rect -10600 -1480 -10560 -1400
rect -10600 -1520 -10300 -1480
rect 5700 -1520 5800 -1480
rect -10600 -1600 -10560 -1520
rect -10600 -1640 -10300 -1600
rect 5700 -1640 5800 -1600
rect -10600 -1720 -10560 -1640
rect -10600 -1760 -10300 -1720
rect 5700 -1760 5800 -1720
rect -10600 -1840 -10560 -1760
rect -10600 -1880 -10300 -1840
rect 5700 -1880 5800 -1840
rect -10600 -1960 -10560 -1880
rect -10600 -2000 -10300 -1960
rect 5700 -2000 5800 -1960
rect -10600 -2080 -10560 -2000
rect -10600 -2120 -10300 -2080
rect 5700 -2120 5800 -2080
rect -10600 -2200 -10560 -2120
rect -10600 -2240 -10300 -2200
rect 5700 -2240 5800 -2200
rect -10600 -2320 -10560 -2240
rect -10600 -2360 -10300 -2320
rect 5700 -2360 5800 -2320
rect -10600 -2440 -10560 -2360
rect -10600 -2480 -10300 -2440
rect 5700 -2480 5800 -2440
rect -10600 -2560 -10560 -2480
rect -10600 -2600 -10300 -2560
rect 5700 -2600 5800 -2560
rect -10600 -2680 -10560 -2600
rect -10600 -2720 -10300 -2680
rect 5700 -2720 5800 -2680
rect -10600 -2800 -10560 -2720
rect -10600 -2840 -10300 -2800
rect 5700 -2840 5800 -2800
rect -10600 -2920 -10560 -2840
rect -10600 -2960 -10300 -2920
rect 5700 -2960 5800 -2920
rect -10600 -3040 -10560 -2960
rect -10600 -3080 -10300 -3040
rect 5700 -3080 5800 -3040
rect -10600 -3160 -10560 -3080
rect -10600 -3200 -10300 -3160
rect 5700 -3200 5800 -3160
rect -10600 -3280 -10560 -3200
rect -10600 -3320 -10300 -3280
rect 5700 -3320 5800 -3280
rect -10600 -3400 -10560 -3320
rect -10600 -3440 -10300 -3400
rect 5700 -3440 5800 -3400
rect -10600 -3520 -10560 -3440
rect -10600 -3560 -10300 -3520
rect 5700 -3560 5800 -3520
rect -10600 -3640 -10560 -3560
rect -10600 -3680 -10300 -3640
rect 5700 -3680 5800 -3640
rect -10600 -3760 -10560 -3680
rect -10600 -3800 -10300 -3760
rect 5700 -3800 5800 -3760
rect -10600 -3880 -10560 -3800
rect -10600 -3920 -10300 -3880
rect 5700 -3920 5800 -3880
rect -10600 -4000 -10560 -3920
rect -10600 -4040 -10300 -4000
rect 5700 -4040 5800 -4000
rect -10600 -4120 -10560 -4040
rect -10600 -4160 -10300 -4120
rect 5700 -4160 5800 -4120
rect -10600 -4240 -10560 -4160
rect -10600 -4280 -10300 -4240
rect 5700 -4280 5800 -4240
rect -10600 -4360 -10560 -4280
rect -10600 -4400 -10300 -4360
rect 5700 -4400 5800 -4360
rect -10600 -4480 -10560 -4400
rect -10600 -4520 -10300 -4480
rect 5700 -4520 5800 -4480
rect -10600 -4600 -10560 -4520
rect -10600 -4640 -10300 -4600
rect 5700 -4640 5800 -4600
rect -10600 -4720 -10560 -4640
rect -10600 -4760 -10300 -4720
rect 5700 -4760 5800 -4720
rect -10600 -4840 -10560 -4760
rect -10600 -4880 -10300 -4840
rect 5700 -4880 5800 -4840
rect -10600 -4960 -10560 -4880
rect -10600 -5000 -10300 -4960
rect 5700 -5000 5800 -4960
rect -10600 -5080 -10560 -5000
rect -10600 -5120 -10300 -5080
rect 5700 -5120 5800 -5080
rect -10600 -5200 -10560 -5120
rect -10600 -5240 -10300 -5200
rect 5700 -5240 5800 -5200
rect -10600 -5320 -10560 -5240
rect -10600 -5360 -10300 -5320
rect 5700 -5360 5800 -5320
rect -10600 -5440 -10560 -5360
rect -10600 -5480 -10300 -5440
rect 5700 -5480 5800 -5440
rect -10600 -5560 -10560 -5480
rect -10600 -5600 -10300 -5560
rect 5700 -5600 5800 -5560
rect -10600 -5680 -10560 -5600
rect -10600 -5720 -10300 -5680
rect 5700 -5720 5800 -5680
rect -10600 -5800 -10560 -5720
rect -10600 -5840 -10300 -5800
rect 5700 -5840 5800 -5800
rect -10600 -5920 -10560 -5840
rect -10600 -5960 -10300 -5920
rect 5700 -5960 5800 -5920
rect -10600 -6040 -10560 -5960
rect -10600 -6080 -10300 -6040
rect 5700 -6080 5800 -6040
rect -10600 -6160 -10560 -6080
rect -10600 -6200 -10300 -6160
rect 5700 -6200 5800 -6160
rect -10600 -6280 -10560 -6200
rect -10600 -6320 -10300 -6280
rect 5700 -6320 5800 -6280
rect -10600 -6400 -10560 -6320
rect -10600 -6440 -10300 -6400
rect 5700 -6440 5800 -6400
rect -10600 -6520 -10560 -6440
rect -10600 -6560 -10300 -6520
rect 5700 -6560 5800 -6520
rect -10600 -6640 -10560 -6560
rect -10600 -6680 -10300 -6640
rect 5700 -6680 5800 -6640
rect -10600 -6760 -10560 -6680
rect -10600 -6800 -10300 -6760
rect 5700 -6800 5800 -6760
rect -10600 -6880 -10560 -6800
rect -10600 -6920 -10300 -6880
rect 5700 -6920 5800 -6880
rect -10600 -7000 -10560 -6920
rect -10600 -7040 -10300 -7000
rect 5700 -7040 5800 -7000
rect -10600 -7120 -10560 -7040
rect -10600 -7160 -10300 -7120
rect 5700 -7160 5800 -7120
rect -10600 -7240 -10560 -7160
rect -10600 -7280 -10300 -7240
rect 5700 -7280 5800 -7240
rect -10600 -7360 -10560 -7280
rect -10600 -7400 -10300 -7360
rect 5700 -7400 5800 -7360
rect -10600 -7480 -10560 -7400
rect -10600 -7520 -10300 -7480
rect 5700 -7520 5800 -7480
rect -10600 -7600 -10560 -7520
rect -10600 -7640 -10300 -7600
rect 5700 -7640 5800 -7600
rect -10600 -7720 -10560 -7640
rect -10600 -7760 -10300 -7720
rect 5700 -7760 5800 -7720
rect -10600 -7840 -10560 -7760
rect -10600 -7880 -10300 -7840
rect 5700 -7880 5800 -7840
rect -10600 -7960 -10560 -7880
rect -10600 -8000 -10300 -7960
rect 5700 -8000 5800 -7960
rect -10600 -8080 -10560 -8000
rect -10600 -8120 -10300 -8080
rect 5700 -8120 5800 -8080
rect -10600 -8200 -10560 -8120
rect -10600 -8240 -10300 -8200
rect 5700 -8240 5800 -8200
rect -10600 -8320 -10560 -8240
rect -10600 -8360 -10300 -8320
rect 5700 -8360 5800 -8320
rect -10600 -8440 -10560 -8360
rect -10600 -8480 -10300 -8440
rect 5700 -8480 5800 -8440
rect -10600 -8560 -10560 -8480
rect -10600 -8600 -10300 -8560
rect 5700 -8600 5800 -8560
rect -10600 -8680 -10560 -8600
rect -10600 -8720 -10300 -8680
rect 5700 -8720 5800 -8680
rect -10600 -8800 -10560 -8720
rect -10600 -8840 -10300 -8800
rect 5700 -8840 5800 -8800
rect -10600 -8920 -10560 -8840
rect -10600 -8960 -10300 -8920
rect 5700 -8960 5800 -8920
rect -10600 -9040 -10560 -8960
rect -10600 -9080 -10300 -9040
rect 5700 -9080 5800 -9040
rect -10600 -9160 -10560 -9080
rect -10600 -9200 -10300 -9160
rect 5700 -9200 5800 -9160
rect -10600 -9280 -10560 -9200
rect -10600 -9320 -10300 -9280
rect 5700 -9320 5800 -9280
rect -10600 -9400 -10560 -9320
rect -10600 -9440 -10300 -9400
rect 5700 -9440 5800 -9400
rect -10600 -9520 -10560 -9440
rect -10600 -9560 -10300 -9520
rect 5700 -9560 5800 -9520
rect -10600 -9640 -10560 -9560
rect -10600 -9680 -10300 -9640
rect 5700 -9680 5800 -9640
rect -10600 -9760 -10560 -9680
rect -10680 -9800 -10300 -9760
rect 5700 -9800 5800 -9760
<< polycont >>
rect -10640 -9760 -10600 -320
<< locali >>
rect -10480 -220 5700 -200
rect -10480 -260 -10280 -220
rect 5680 -260 5700 -220
rect -10480 -280 5700 -260
rect -10680 -320 -10560 -280
rect -10680 -9760 -10640 -320
rect -10600 -9760 -10560 -320
rect -10680 -9800 -10560 -9760
rect -10480 -440 -10400 -280
rect -10300 -340 5920 -320
rect -10300 -380 -10280 -340
rect 5680 -380 5920 -340
rect -10300 -400 5920 -380
rect -10480 -460 5700 -440
rect -10480 -500 -10280 -460
rect 5680 -500 5700 -460
rect -10480 -520 5700 -500
rect -10480 -680 -10400 -520
rect 5800 -560 5920 -400
rect -10300 -580 5920 -560
rect -10300 -620 -10280 -580
rect 5680 -620 5920 -580
rect -10300 -640 5920 -620
rect -10480 -700 5700 -680
rect -10480 -740 -10280 -700
rect 5680 -740 5700 -700
rect -10480 -760 5700 -740
rect -10480 -920 -10400 -760
rect 5800 -800 5920 -640
rect -10300 -820 5920 -800
rect -10300 -860 -10280 -820
rect 5680 -860 5920 -820
rect -10300 -880 5920 -860
rect -10480 -940 5700 -920
rect -10480 -980 -10280 -940
rect 5680 -980 5700 -940
rect -10480 -1000 5700 -980
rect -10480 -1160 -10400 -1000
rect 5800 -1040 5920 -880
rect -10300 -1060 5920 -1040
rect -10300 -1100 -10280 -1060
rect 5680 -1100 5920 -1060
rect -10300 -1120 5920 -1100
rect -10480 -1180 5700 -1160
rect -10480 -1220 -10280 -1180
rect 5680 -1220 5700 -1180
rect -10480 -1240 5700 -1220
rect -10480 -1400 -10400 -1240
rect 5800 -1280 5920 -1120
rect -10300 -1300 5920 -1280
rect -10300 -1340 -10280 -1300
rect 5680 -1340 5920 -1300
rect -10300 -1360 5920 -1340
rect -10480 -1420 5700 -1400
rect -10480 -1460 -10280 -1420
rect 5680 -1460 5700 -1420
rect -10480 -1480 5700 -1460
rect -10480 -1640 -10400 -1480
rect 5800 -1520 5920 -1360
rect -10300 -1540 5920 -1520
rect -10300 -1580 -10280 -1540
rect 5680 -1580 5920 -1540
rect -10300 -1600 5920 -1580
rect -10480 -1660 5700 -1640
rect -10480 -1700 -10280 -1660
rect 5680 -1700 5700 -1660
rect -10480 -1720 5700 -1700
rect -10480 -1880 -10400 -1720
rect 5800 -1760 5920 -1600
rect -10300 -1780 5920 -1760
rect -10300 -1820 -10280 -1780
rect 5680 -1820 5920 -1780
rect -10300 -1840 5920 -1820
rect -10480 -1900 5700 -1880
rect -10480 -1940 -10280 -1900
rect 5680 -1940 5700 -1900
rect -10480 -1960 5700 -1940
rect -10480 -2120 -10400 -1960
rect 5800 -2000 5920 -1840
rect -10300 -2020 5920 -2000
rect -10300 -2060 -10280 -2020
rect 5680 -2060 5920 -2020
rect -10300 -2080 5920 -2060
rect -10480 -2140 5700 -2120
rect -10480 -2180 -10280 -2140
rect 5680 -2180 5700 -2140
rect -10480 -2200 5700 -2180
rect -10480 -2360 -10400 -2200
rect 5800 -2240 5920 -2080
rect -10300 -2260 5920 -2240
rect -10300 -2300 -10280 -2260
rect 5680 -2300 5920 -2260
rect -10300 -2320 5920 -2300
rect -10480 -2380 5700 -2360
rect -10480 -2420 -10280 -2380
rect 5680 -2420 5700 -2380
rect -10480 -2440 5700 -2420
rect -10480 -2600 -10400 -2440
rect 5800 -2480 5920 -2320
rect -10300 -2500 5920 -2480
rect -10300 -2540 -10280 -2500
rect 5680 -2540 5920 -2500
rect -10300 -2560 5920 -2540
rect -10480 -2620 5700 -2600
rect -10480 -2660 -10280 -2620
rect 5680 -2660 5700 -2620
rect -10480 -2680 5700 -2660
rect -10480 -2840 -10400 -2680
rect 5800 -2720 5920 -2560
rect -10300 -2740 5920 -2720
rect -10300 -2780 -10280 -2740
rect 5680 -2780 5920 -2740
rect -10300 -2800 5920 -2780
rect -10480 -2860 5700 -2840
rect -10480 -2900 -10280 -2860
rect 5680 -2900 5700 -2860
rect -10480 -2920 5700 -2900
rect -10480 -3080 -10400 -2920
rect 5800 -2960 5920 -2800
rect -10300 -2980 5920 -2960
rect -10300 -3020 -10280 -2980
rect 5680 -3020 5920 -2980
rect -10300 -3040 5920 -3020
rect -10480 -3100 5700 -3080
rect -10480 -3140 -10280 -3100
rect 5680 -3140 5700 -3100
rect -10480 -3160 5700 -3140
rect -10480 -3320 -10400 -3160
rect 5800 -3200 5920 -3040
rect -10300 -3220 5920 -3200
rect -10300 -3260 -10280 -3220
rect 5680 -3260 5920 -3220
rect -10300 -3280 5920 -3260
rect -10480 -3340 5700 -3320
rect -10480 -3380 -10280 -3340
rect 5680 -3380 5700 -3340
rect -10480 -3400 5700 -3380
rect -10480 -3560 -10400 -3400
rect 5800 -3440 5920 -3280
rect -10300 -3460 5920 -3440
rect -10300 -3500 -10280 -3460
rect 5680 -3500 5920 -3460
rect -10300 -3520 5920 -3500
rect -10480 -3580 5700 -3560
rect -10480 -3620 -10280 -3580
rect 5680 -3620 5700 -3580
rect -10480 -3640 5700 -3620
rect -10480 -3800 -10400 -3640
rect 5800 -3680 5920 -3520
rect -10300 -3700 5920 -3680
rect -10300 -3740 -10280 -3700
rect 5680 -3740 5920 -3700
rect -10300 -3760 5920 -3740
rect -10480 -3820 5700 -3800
rect -10480 -3860 -10280 -3820
rect 5680 -3860 5700 -3820
rect -10480 -3880 5700 -3860
rect -10480 -4040 -10400 -3880
rect 5800 -3920 5920 -3760
rect -10300 -3940 5920 -3920
rect -10300 -3980 -10280 -3940
rect 5680 -3980 5920 -3940
rect -10300 -4000 5920 -3980
rect -10480 -4060 5700 -4040
rect -10480 -4100 -10280 -4060
rect 5680 -4100 5700 -4060
rect -10480 -4120 5700 -4100
rect -10480 -4280 -10400 -4120
rect 5800 -4160 5920 -4000
rect -10300 -4180 5920 -4160
rect -10300 -4220 -10280 -4180
rect 5680 -4220 5920 -4180
rect -10300 -4240 5920 -4220
rect -10480 -4300 5700 -4280
rect -10480 -4340 -10280 -4300
rect 5680 -4340 5700 -4300
rect -10480 -4360 5700 -4340
rect -10480 -4520 -10400 -4360
rect 5800 -4400 5920 -4240
rect -10300 -4420 5920 -4400
rect -10300 -4460 -10280 -4420
rect 5680 -4460 5920 -4420
rect -10300 -4480 5920 -4460
rect -10480 -4540 5700 -4520
rect -10480 -4580 -10280 -4540
rect 5680 -4580 5700 -4540
rect -10480 -4600 5700 -4580
rect -10480 -4760 -10400 -4600
rect 5800 -4640 5920 -4480
rect -10300 -4660 5920 -4640
rect -10300 -4700 -10280 -4660
rect 5680 -4700 5920 -4660
rect -10300 -4720 5920 -4700
rect -10480 -4780 5700 -4760
rect -10480 -4820 -10280 -4780
rect 5680 -4820 5700 -4780
rect -10480 -4840 5700 -4820
rect -10480 -5000 -10400 -4840
rect 5800 -4880 5920 -4720
rect -10300 -4900 5920 -4880
rect -10300 -4940 -10280 -4900
rect 5680 -4940 5920 -4900
rect -10300 -4960 5920 -4940
rect -10480 -5020 5700 -5000
rect -10480 -5060 -10280 -5020
rect 5680 -5060 5700 -5020
rect -10480 -5080 5700 -5060
rect -10480 -5240 -10400 -5080
rect 5800 -5120 5920 -4960
rect -10300 -5140 5920 -5120
rect -10300 -5180 -10280 -5140
rect 5680 -5180 5920 -5140
rect -10300 -5200 5920 -5180
rect -10480 -5260 5700 -5240
rect -10480 -5300 -10280 -5260
rect 5680 -5300 5700 -5260
rect -10480 -5320 5700 -5300
rect -10480 -5480 -10400 -5320
rect 5800 -5360 5920 -5200
rect -10300 -5380 5920 -5360
rect -10300 -5420 -10280 -5380
rect 5680 -5420 5920 -5380
rect -10300 -5440 5920 -5420
rect -10480 -5500 5700 -5480
rect -10480 -5540 -10280 -5500
rect 5680 -5540 5700 -5500
rect -10480 -5560 5700 -5540
rect -10480 -5720 -10400 -5560
rect 5800 -5600 5920 -5440
rect -10300 -5620 5920 -5600
rect -10300 -5660 -10280 -5620
rect 5680 -5660 5920 -5620
rect -10300 -5680 5920 -5660
rect -10480 -5740 5700 -5720
rect -10480 -5780 -10280 -5740
rect 5680 -5780 5700 -5740
rect -10480 -5800 5700 -5780
rect -10480 -5960 -10400 -5800
rect 5800 -5840 5920 -5680
rect -10300 -5860 5920 -5840
rect -10300 -5900 -10280 -5860
rect 5680 -5900 5920 -5860
rect -10300 -5920 5920 -5900
rect -10480 -5980 5700 -5960
rect -10480 -6020 -10280 -5980
rect 5680 -6020 5700 -5980
rect -10480 -6040 5700 -6020
rect -10480 -6200 -10400 -6040
rect 5800 -6080 5920 -5920
rect -10300 -6100 5920 -6080
rect -10300 -6140 -10280 -6100
rect 5680 -6140 5920 -6100
rect -10300 -6160 5920 -6140
rect -10480 -6220 5700 -6200
rect -10480 -6260 -10280 -6220
rect 5680 -6260 5700 -6220
rect -10480 -6280 5700 -6260
rect -10480 -6440 -10400 -6280
rect 5800 -6320 5920 -6160
rect -10300 -6340 5920 -6320
rect -10300 -6380 -10280 -6340
rect 5680 -6380 5920 -6340
rect -10300 -6400 5920 -6380
rect -10480 -6460 5700 -6440
rect -10480 -6500 -10280 -6460
rect 5680 -6500 5700 -6460
rect -10480 -6520 5700 -6500
rect -10480 -6680 -10400 -6520
rect 5800 -6560 5920 -6400
rect -10300 -6580 5920 -6560
rect -10300 -6620 -10280 -6580
rect 5680 -6620 5920 -6580
rect -10300 -6640 5920 -6620
rect -10480 -6700 5700 -6680
rect -10480 -6740 -10280 -6700
rect 5680 -6740 5700 -6700
rect -10480 -6760 5700 -6740
rect -10480 -6920 -10400 -6760
rect 5800 -6800 5920 -6640
rect -10300 -6820 5920 -6800
rect -10300 -6860 -10280 -6820
rect 5680 -6860 5920 -6820
rect -10300 -6880 5920 -6860
rect -10480 -6940 5700 -6920
rect -10480 -6980 -10280 -6940
rect 5680 -6980 5700 -6940
rect -10480 -7000 5700 -6980
rect -10480 -7160 -10400 -7000
rect 5800 -7040 5920 -6880
rect -10300 -7060 5920 -7040
rect -10300 -7100 -10280 -7060
rect 5680 -7100 5920 -7060
rect -10300 -7120 5920 -7100
rect -10480 -7180 5700 -7160
rect -10480 -7220 -10280 -7180
rect 5680 -7220 5700 -7180
rect -10480 -7240 5700 -7220
rect -10480 -7400 -10400 -7240
rect 5800 -7280 5920 -7120
rect -10300 -7300 5920 -7280
rect -10300 -7340 -10280 -7300
rect 5680 -7340 5920 -7300
rect -10300 -7360 5920 -7340
rect -10480 -7420 5700 -7400
rect -10480 -7460 -10280 -7420
rect 5680 -7460 5700 -7420
rect -10480 -7480 5700 -7460
rect -10480 -7640 -10400 -7480
rect 5800 -7520 5920 -7360
rect -10300 -7540 5920 -7520
rect -10300 -7580 -10280 -7540
rect 5680 -7580 5920 -7540
rect -10300 -7600 5920 -7580
rect -10480 -7660 5700 -7640
rect -10480 -7700 -10280 -7660
rect 5680 -7700 5700 -7660
rect -10480 -7720 5700 -7700
rect -10480 -7880 -10400 -7720
rect 5800 -7760 5920 -7600
rect -10300 -7780 5920 -7760
rect -10300 -7820 -10280 -7780
rect 5680 -7820 5920 -7780
rect -10300 -7840 5920 -7820
rect -10480 -7900 5700 -7880
rect -10480 -7940 -10280 -7900
rect 5680 -7940 5700 -7900
rect -10480 -7960 5700 -7940
rect -10480 -8120 -10400 -7960
rect 5800 -8000 5920 -7840
rect -10300 -8020 5920 -8000
rect -10300 -8060 -10280 -8020
rect 5680 -8060 5920 -8020
rect -10300 -8080 5920 -8060
rect -10480 -8140 5700 -8120
rect -10480 -8180 -10280 -8140
rect 5680 -8180 5700 -8140
rect -10480 -8200 5700 -8180
rect -10480 -8360 -10400 -8200
rect 5800 -8240 5920 -8080
rect -10300 -8260 5920 -8240
rect -10300 -8300 -10280 -8260
rect 5680 -8300 5920 -8260
rect -10300 -8320 5920 -8300
rect -10480 -8380 5700 -8360
rect -10480 -8420 -10280 -8380
rect 5680 -8420 5700 -8380
rect -10480 -8440 5700 -8420
rect -10480 -8600 -10400 -8440
rect 5800 -8480 5920 -8320
rect -10300 -8500 5920 -8480
rect -10300 -8540 -10280 -8500
rect 5680 -8540 5920 -8500
rect -10300 -8560 5920 -8540
rect -10480 -8620 5700 -8600
rect -10480 -8660 -10280 -8620
rect 5680 -8660 5700 -8620
rect -10480 -8680 5700 -8660
rect -10480 -8840 -10400 -8680
rect 5800 -8720 5920 -8560
rect -10300 -8740 5920 -8720
rect -10300 -8780 -10280 -8740
rect 5680 -8780 5920 -8740
rect -10300 -8800 5920 -8780
rect -10480 -8860 5700 -8840
rect -10480 -8900 -10280 -8860
rect 5680 -8900 5700 -8860
rect -10480 -8920 5700 -8900
rect -10480 -9080 -10400 -8920
rect 5800 -8960 5920 -8800
rect -10300 -8980 5920 -8960
rect -10300 -9020 -10280 -8980
rect 5680 -9020 5920 -8980
rect -10300 -9040 5920 -9020
rect -10480 -9100 5700 -9080
rect -10480 -9140 -10280 -9100
rect 5680 -9140 5700 -9100
rect -10480 -9160 5700 -9140
rect -10480 -9320 -10400 -9160
rect 5800 -9200 5920 -9040
rect -10300 -9220 5920 -9200
rect -10300 -9260 -10280 -9220
rect 5680 -9260 5920 -9220
rect -10300 -9280 5920 -9260
rect -10480 -9340 5700 -9320
rect -10480 -9380 -10280 -9340
rect 5680 -9380 5700 -9340
rect -10480 -9400 5700 -9380
rect -10480 -9560 -10400 -9400
rect 5800 -9440 5920 -9280
rect -10300 -9460 5920 -9440
rect -10300 -9500 -10280 -9460
rect 5680 -9500 5920 -9460
rect -10300 -9520 5920 -9500
rect -10480 -9580 5700 -9560
rect -10480 -9620 -10280 -9580
rect 5680 -9620 5700 -9580
rect -10480 -9640 5700 -9620
rect -10480 -9800 -10400 -9640
rect 5800 -9680 5920 -9520
rect -10300 -9700 5920 -9680
rect -10300 -9740 -10280 -9700
rect 5680 -9740 5920 -9700
rect -10300 -9760 5920 -9740
rect -10480 -9820 5700 -9800
rect -10480 -9860 -10280 -9820
rect 5680 -9860 5700 -9820
rect -10480 -9880 5700 -9860
<< labels >>
flabel pdiffc -3120 -240 -3120 -240 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont -10625 -3478 -10625 -3478 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel locali 5859 -5501 5859 -5501 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel nwell -10717 -200 -10717 -200 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
