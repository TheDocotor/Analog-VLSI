magic
tech sky130A
magscale 1 2
timestamp 1732122809
<< nwell >>
rect -894 -598 894 564
<< pmos >>
rect -800 -536 800 464
<< pdiff >>
rect -858 452 -800 464
rect -858 -524 -846 452
rect -812 -524 -800 452
rect -858 -536 -800 -524
rect 800 452 858 464
rect 800 -524 812 452
rect 846 -524 858 452
rect 800 -536 858 -524
<< pdiffc >>
rect -846 -524 -812 452
rect 812 -524 846 452
<< poly >>
rect -800 545 800 561
rect -800 511 -784 545
rect 784 511 800 545
rect -800 464 800 511
rect -800 -562 800 -536
<< polycont >>
rect -784 511 784 545
<< locali >>
rect -800 511 -784 545
rect 784 511 800 545
rect -846 452 -812 468
rect -846 -540 -812 -524
rect 812 452 846 468
rect 812 -540 846 -524
<< viali >>
rect -784 511 784 545
rect -846 -524 -812 452
rect 812 -524 846 452
<< metal1 >>
rect -796 545 796 551
rect -796 511 -784 545
rect 784 511 796 545
rect -796 505 796 511
rect -852 452 -806 464
rect -852 -524 -846 452
rect -812 -524 -806 452
rect -852 -536 -806 -524
rect 806 452 852 464
rect 806 -524 812 452
rect 846 -524 852 452
rect 806 -536 852 -524
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_01v8_GXDZBM parameters
<< end >>
