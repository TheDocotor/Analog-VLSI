magic
tech sky130A
magscale 1 2
timestamp 1733333627
<< locali >>
rect -2400 17520 -1600 27500
rect -2400 17440 21740 17520
rect -2400 1800 -1600 17440
<< viali >>
rect 1800 32000 2200 32200
rect 5240 28720 5440 28820
rect 7550 28750 7670 28810
rect -7406 25618 -6726 25858
rect -11000 25000 -10600 25200
rect 3534 26446 3702 26480
rect -500 23600 -300 23900
rect 14800 23400 15100 23600
rect 656 21727 764 22127
rect 956 21727 1064 22127
rect 7500 18560 7540 19540
rect 1280 18260 1410 18370
rect 7440 16880 7580 16980
rect 14700 16000 15000 16200
<< metal1 >>
rect -22200 26200 -21400 26600
rect -17900 25200 -9800 25500
rect 2600 25480 2900 25660
rect -17900 25000 -11000 25200
rect -10600 25000 -9800 25200
rect -17900 24900 -9800 25000
rect -44 22127 62 22535
rect 256 22127 362 22535
rect 20820 19840 20900 20040
rect 7460 19520 7500 19540
rect 7460 18560 7480 19520
rect 7540 18560 7560 19540
rect 7460 18520 7560 18560
rect -1240 13660 -1120 14040
rect 24800 12440 24940 12640
rect 25480 11792 25718 12014
<< via1 >>
rect 1800 32000 2200 32200
rect 5240 28720 5440 28820
rect 7550 28750 7670 28810
rect 3534 26446 3702 26480
rect -7406 25618 -6726 25858
rect -11000 25000 -10600 25200
rect -500 23600 -300 23900
rect 14800 23400 15100 23600
rect 656 21727 764 22127
rect 956 21727 1064 22127
rect 7480 18560 7500 19520
rect 7500 18560 7540 19520
rect 1280 18260 1410 18370
rect 7440 16880 7580 16980
rect 14700 16000 15000 16200
<< metal2 >>
rect 1700 32200 2300 32300
rect -3600 32000 1800 32200
rect 2200 32000 2300 32200
rect -3600 27800 -3400 32000
rect 1700 31900 2300 32000
rect 7530 28810 7690 28830
rect 7530 28750 7550 28810
rect 7670 28750 7690 28810
rect 7530 28730 7690 28750
rect -11000 27600 -3400 27800
rect -11000 25300 -10600 27600
rect 3600 26480 3700 26500
rect 3600 26300 3700 26446
rect -7200 26200 3700 26300
rect -7200 25858 -6800 26200
rect -7200 25600 -6800 25618
rect -11100 25200 -10500 25300
rect -11100 25000 -11000 25200
rect -10600 25000 -10500 25200
rect -11100 24900 -10500 25000
rect -5600 18400 -5100 26200
rect -600 23900 -200 24000
rect -600 23600 -500 23900
rect -300 23600 -200 23900
rect -600 23500 -200 23600
rect 14700 23600 15200 23700
rect 14700 23400 14800 23600
rect 15100 23400 15200 23600
rect 14700 23300 15200 23400
rect 7460 19520 7560 19540
rect 7460 18560 7480 19520
rect 7540 18560 7560 19520
rect 7460 18520 7560 18560
rect -5600 18370 1400 18400
rect -5600 18260 1280 18370
rect -5600 18200 1400 18260
rect 7420 16980 7600 17000
rect 7420 16880 7440 16980
rect 7580 16880 7600 16980
rect 7420 16860 7600 16880
rect 14600 16200 15100 16300
rect 14600 16000 14700 16200
rect 15000 16000 15100 16200
rect 14600 15900 15100 16000
<< via2 >>
rect 5240 28720 5440 28820
rect 7550 28750 7670 28810
rect -11000 25000 -10600 25200
rect -500 23600 -300 23900
rect 14800 23400 15100 23600
rect 656 21727 764 22127
rect 956 21727 1064 22127
rect 7480 18560 7540 19520
rect 7440 16880 7580 16980
rect 14700 16000 15000 16200
<< metal3 >>
rect 5220 28820 5460 28840
rect 5220 28800 5240 28820
rect 5200 28720 5240 28800
rect 5440 28720 5460 28820
rect 7520 28810 7680 28820
rect 7520 28800 7550 28810
rect 5200 28700 5460 28720
rect 7500 28750 7550 28800
rect 7670 28800 7680 28810
rect 7670 28750 7700 28800
rect -11100 25200 -1700 25300
rect -11100 25000 -11000 25200
rect -10600 25000 -1700 25200
rect -11100 24900 -1700 25000
rect -2100 24000 -1700 24900
rect -2100 23900 -200 24000
rect 5200 23900 5400 28700
rect -2100 23600 -500 23900
rect -300 23600 -200 23900
rect -2100 23500 -200 23600
rect 900 23600 5400 23900
rect 600 22127 800 22200
rect 600 21727 656 22127
rect 764 21727 800 22127
rect 600 21600 800 21727
rect 900 22127 1100 23600
rect 7500 23400 7700 28750
rect 900 21727 956 22127
rect 1064 21727 1100 22127
rect 900 21700 1100 21727
rect 1500 23200 7700 23400
rect 14600 23600 15200 23700
rect 14600 23400 14800 23600
rect 15100 23400 15200 23600
rect 1500 21600 1700 23200
rect 600 21400 1700 21600
rect 7460 19520 7560 19540
rect 7460 18560 7480 19520
rect 7540 18560 7560 19520
rect 7460 18520 7560 18560
rect 7460 17000 7540 18520
rect 7420 16980 7600 17000
rect 7420 16880 7440 16980
rect 7580 16880 7600 16980
rect 7420 16860 7600 16880
rect 14600 16200 15200 23400
rect 14600 16000 14700 16200
rect 15000 16000 15200 16200
rect 14600 15900 15200 16000
use bandgap  bandgap_0 ~/Documents/ece5120/hw05/mag
timestamp 1732920865
transform 1 0 -15746 0 1 19418
box -6800 -18000 13400 8100
use demod  demod_0 ~/Documents/ece5120/hw08/mag
timestamp 1733331218
transform 1 0 -5460 0 1 13840
box 1300 -13500 32200 3600
use gill_cell  gill_cell_0 ~/Documents/ece5120/hw07/mag
timestamp 1732920865
transform 1 0 1540 0 1 22520
box -3200 -5000 20200 2400
use lna  lna_0 ~/Documents/ece5120/hw06/mag
timestamp 1733178114
transform 1 0 3940 0 1 26120
box -5600 -1200 18400 6800
<< labels >>
flabel via1 -7060 25720 -7060 25720 0 FreeSans 1600 0 0 0 Vref
port 7 nsew
flabel metal1 20860 19940 20860 19940 0 FreeSans 1600 0 0 0 IF_out
port 3 nsew
flabel metal1 300 22520 300 22520 0 FreeSans 1600 0 0 0 LOp
port 4 nsew
flabel metal1 0 22280 0 22280 0 FreeSans 1600 0 0 0 LOn
port 5 nsew
flabel via2 7500 16940 7500 16940 0 FreeSans 1600 0 0 0 RFn
flabel metal1 -1200 13800 -1200 13800 0 FreeSans 1600 0 0 0 IF_in
port 2 nsew
flabel metal1 2800 25600 2800 25600 0 FreeSans 1600 0 0 0 ANT
port 1 nsew
flabel metal1 -21900 26400 -21900 26400 0 FreeSans 1600 0 0 0 VSS
port 8 nsew
flabel metal1 -14000 25200 -14000 25200 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal1 25598 11912 25598 11912 0 FreeSans 1600 0 0 0 RC
port 9 nsew
<< end >>
