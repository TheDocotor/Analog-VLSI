magic
tech sky130A
magscale 1 2
timestamp 1730763316
<< nwell >>
rect -225 -1150 1075 550
<< pmos >>
rect 100 200 900 400
rect 100 -100 900 100
rect 100 -400 900 -200
rect 100 -700 900 -500
rect 100 -1000 900 -800
<< pdiff >>
rect 100 475 900 500
rect 100 425 125 475
rect 875 425 900 475
rect 100 400 900 425
rect 100 175 900 200
rect 100 125 125 175
rect 875 125 900 175
rect 100 100 900 125
rect 100 -125 900 -100
rect 100 -175 125 -125
rect 875 -175 900 -125
rect 100 -200 900 -175
rect 100 -425 900 -400
rect 100 -475 125 -425
rect 875 -475 900 -425
rect 100 -500 900 -475
rect 100 -725 900 -700
rect 100 -775 125 -725
rect 875 -775 900 -725
rect 100 -800 900 -775
rect 100 -1025 900 -1000
rect 100 -1075 125 -1025
rect 875 -1075 900 -1025
rect 100 -1100 900 -1075
<< pdiffc >>
rect 125 425 875 475
rect 125 125 875 175
rect 125 -175 875 -125
rect 125 -475 875 -425
rect 125 -775 875 -725
rect 125 -1075 875 -1025
<< poly >>
rect -200 375 100 400
rect -200 -975 -175 375
rect -125 200 100 375
rect 900 200 1000 400
rect -125 100 0 200
rect -125 -100 100 100
rect 900 -100 1000 100
rect -125 -200 0 -100
rect -125 -400 100 -200
rect 900 -400 1000 -200
rect -125 -500 0 -400
rect -125 -700 100 -500
rect 900 -700 1000 -500
rect -125 -800 0 -700
rect -125 -975 100 -800
rect -200 -1000 100 -975
rect 900 -1000 1000 -800
<< polycont >>
rect -175 -975 -125 375
<< locali >>
rect -50 475 900 500
rect -50 425 125 475
rect 875 425 900 475
rect -50 400 900 425
rect -200 375 -100 400
rect -200 -975 -175 375
rect -125 -975 -100 375
rect -50 -100 50 400
rect 100 175 1050 200
rect 100 125 125 175
rect 875 125 1050 175
rect 100 100 1050 125
rect -50 -125 900 -100
rect -50 -175 125 -125
rect 875 -175 900 -125
rect -50 -200 900 -175
rect -50 -700 50 -200
rect 950 -400 1050 100
rect 100 -425 1050 -400
rect 100 -475 125 -425
rect 875 -475 1050 -425
rect 100 -500 1050 -475
rect -50 -725 900 -700
rect -50 -775 125 -725
rect 875 -775 900 -725
rect -50 -800 900 -775
rect -200 -1000 -100 -975
rect 950 -1000 1050 -500
rect 100 -1025 1050 -1000
rect 100 -1075 125 -1025
rect 875 -1075 1050 -1025
rect 100 -1100 1050 -1075
<< labels >>
flabel pdiffc 600 450 600 450 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel pdiffc 625 -1050 625 -1050 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel polycont -150 -300 -150 -300 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel nwell -150 475 -150 475 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
