magic
tech sky130A
magscale 1 2
timestamp 1730254111
<< nwell >>
rect -100 -1100 1200 700
<< pmos >>
rect 100 300 1000 500
rect 100 0 1000 200
rect 100 -300 1000 -100
rect 100 -600 1000 -400
rect 100 -900 1000 -700
<< pdiff >>
rect 100 575 1000 600
rect 100 525 125 575
rect 975 525 1000 575
rect 100 500 1000 525
rect 100 275 1000 300
rect 100 225 125 275
rect 975 225 1000 275
rect 100 200 1000 225
rect 100 -25 1000 0
rect 100 -75 125 -25
rect 975 -75 1000 -25
rect 100 -100 1000 -75
rect 100 -325 1000 -300
rect 100 -375 125 -325
rect 975 -375 1000 -325
rect 100 -400 1000 -375
rect 100 -625 1000 -600
rect 100 -675 125 -625
rect 975 -675 1000 -625
rect 100 -700 1000 -675
rect 100 -925 1000 -900
rect 100 -975 125 -925
rect 975 -975 1000 -925
rect 100 -1000 1000 -975
<< pdiffc >>
rect 125 525 975 575
rect 125 225 975 275
rect 125 -75 975 -25
rect 125 -375 975 -325
rect 125 -675 975 -625
rect 125 -975 975 -925
<< poly >>
rect 0 300 100 500
rect 1000 300 1100 500
rect 0 0 100 200
rect 1000 0 1100 200
rect 0 -300 100 -100
rect 1000 -300 1100 -100
rect 0 -600 100 -400
rect 1000 -600 1100 -400
rect 0 -900 100 -700
rect 1000 -900 1100 -700
<< locali >>
rect 100 575 1000 600
rect 100 525 125 575
rect 975 525 1000 575
rect 100 500 1000 525
rect 100 275 1000 300
rect 100 225 125 275
rect 975 225 1000 275
rect 100 200 1000 225
rect 100 -25 1000 0
rect 100 -75 125 -25
rect 975 -75 1000 -25
rect 100 -100 1000 -75
rect 100 -325 1000 -300
rect 100 -375 125 -325
rect 975 -375 1000 -325
rect 100 -400 1000 -375
rect 100 -625 1000 -600
rect 100 -675 125 -625
rect 975 -675 1000 -625
rect 100 -700 1000 -675
rect 100 -925 1000 -900
rect 100 -975 125 -925
rect 975 -975 1000 -925
rect 100 -1000 1000 -975
<< end >>
