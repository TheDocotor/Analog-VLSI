magic
tech sky130A
magscale 1 2
timestamp 1731518900
<< nwell >>
rect -1400 -1200 3200 1000
<< nsubdiff >>
rect -1350 800 0 900
rect 1700 800 3150 900
rect -1350 550 -1250 800
rect -1350 -1050 -1250 -900
rect 3050 500 3150 800
rect 3050 -1050 3150 -850
rect -1350 -1150 100 -1050
rect 1900 -1150 3150 -1050
<< nsubdiffcont >>
rect 0 800 1700 900
rect -1350 -900 -1250 550
rect 3050 -850 3150 500
rect 100 -1150 1900 -1050
<< locali >>
rect -1350 800 0 900
rect 1700 800 3150 900
rect -1350 550 -1250 800
rect 700 550 1050 650
rect -1350 -1050 -1250 -900
rect 3050 500 3150 800
rect 3050 -1050 3150 -850
rect -1350 -1150 100 -1050
rect 1900 -1150 3150 -1050
use p40x1  p40x1_0
timestamp 1731517860
transform 1 0 1025 0 1 150
box -225 -1150 1875 550
use p40x1  p40x1_1
timestamp 1731517860
transform -1 0 725 0 1 150
box -225 -1150 1875 550
<< labels >>
flabel nwell 500 600 500 600 0 FreeSans 1600 0 0 0 D
port 0 nsew
flabel nwell 900 -100 900 -100 0 FreeSans 1600 0 0 0 G
port 1 nsew
flabel nwell -150 -900 -150 -900 0 FreeSans 1600 0 0 0 RS
port 2 nsew
flabel nwell 2050 -900 2050 -900 0 FreeSans 1600 0 0 0 LS
port 3 nsew
flabel nwell -1050 850 -1050 850 0 FreeSans 1600 0 0 0 B
port 4 nsew
<< end >>
