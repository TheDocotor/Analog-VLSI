magic
tech sky130A
timestamp 1732735194
<< nwell >>
rect 80 100 690 180
rect 150 -520 410 -420
<< locali >>
rect 80 100 690 180
rect 150 -520 410 -420
use p1x15  p1x15_0
timestamp 1732726409
transform -1 0 -40 0 -1 -320
box -500 -600 500 300
use p1x15  p1x15_1
timestamp 1732726409
transform 1 0 760 0 -1 -320
box -500 -600 500 300
<< labels >>
flabel space -90 -470 -90 -470 0 FreeSans 800 0 0 0 DL
port 1 nsew
flabel space 810 -470 810 -470 0 FreeSans 800 0 0 0 DR
port 2 nsew
flabel space 360 -180 360 -180 0 FreeSans 800 0 0 0 G
port 3 nsew
flabel space -90 130 -90 130 0 FreeSans 800 0 0 0 SL
port 4 nsew
flabel space 820 130 820 130 0 FreeSans 800 0 0 0 SR
port 5 nsew
flabel space -480 200 -480 200 0 FreeSans 800 0 0 0 B
port 6 nsew
<< end >>
