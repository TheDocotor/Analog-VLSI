magic
tech sky130A
magscale 1 2
timestamp 1732757215
<< nmos >>
rect -100 -169 100 231
<< ndiff >>
rect -158 219 -100 231
rect -158 -157 -146 219
rect -112 -157 -100 219
rect -158 -169 -100 -157
rect 100 219 158 231
rect 100 -157 112 219
rect 146 -157 158 219
rect 100 -169 158 -157
<< ndiffc >>
rect -146 -157 -112 219
rect 112 -157 146 219
<< poly >>
rect -100 231 100 257
rect -100 -207 100 -169
rect -100 -241 -84 -207
rect 84 -241 100 -207
rect -100 -257 100 -241
<< polycont >>
rect -84 -241 84 -207
<< locali >>
rect -146 219 -112 235
rect -146 -173 -112 -157
rect 112 219 146 235
rect 112 -173 146 -157
rect -100 -241 -84 -207
rect 84 -241 100 -207
<< viali >>
rect -146 -157 -112 219
rect 112 -157 146 219
rect -84 -241 84 -207
<< metal1 >>
rect -152 219 -106 231
rect -152 -157 -146 219
rect -112 -157 -106 219
rect -152 -169 -106 -157
rect 106 219 152 231
rect 106 -157 112 219
rect 146 -157 152 219
rect 106 -169 152 -157
rect -96 -207 96 -201
rect -96 -241 -84 -207
rect 84 -241 96 -207
rect -96 -247 96 -241
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_Q7B869 parameters
<< end >>
