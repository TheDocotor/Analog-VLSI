magic
tech sky130A
magscale 1 2
timestamp 1732122809
<< nmos >>
rect -200 -531 200 469
<< ndiff >>
rect -258 457 -200 469
rect -258 -519 -246 457
rect -212 -519 -200 457
rect -258 -531 -200 -519
rect 200 457 258 469
rect 200 -519 212 457
rect 246 -519 258 457
rect 200 -531 258 -519
<< ndiffc >>
rect -246 -519 -212 457
rect 212 -519 246 457
<< poly >>
rect -200 541 200 557
rect -200 507 -184 541
rect 184 507 200 541
rect -200 469 200 507
rect -200 -557 200 -531
<< polycont >>
rect -184 507 184 541
<< locali >>
rect -200 507 -184 541
rect 184 507 200 541
rect -246 457 -212 473
rect -246 -535 -212 -519
rect 212 457 246 473
rect 212 -535 246 -519
<< viali >>
rect -184 507 184 541
rect -246 -519 -212 457
rect 212 -519 246 457
<< metal1 >>
rect -196 541 196 547
rect -196 507 -184 541
rect 184 507 196 541
rect -196 501 196 507
rect -252 457 -206 469
rect -252 -519 -246 457
rect -212 -519 -206 457
rect -252 -531 -206 -519
rect 206 457 252 469
rect 206 -519 212 457
rect 246 -519 252 457
rect 206 -531 252 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_8WUFR5 parameters
<< end >>
