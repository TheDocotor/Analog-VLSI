magic
tech sky130A
timestamp 1730605901
<< nmos >>
rect -2500 -21 2500 21
<< ndiff >>
rect -2529 15 -2500 21
rect -2529 -15 -2523 15
rect -2506 -15 -2500 15
rect -2529 -21 -2500 -15
rect 2500 15 2529 21
rect 2500 -15 2506 15
rect 2523 -15 2529 15
rect 2500 -21 2529 -15
<< ndiffc >>
rect -2523 -15 -2506 15
rect 2506 -15 2523 15
<< poly >>
rect -2500 21 2500 34
rect -2500 -34 2500 -21
<< locali >>
rect -2523 15 -2506 23
rect -2523 -23 -2506 -15
rect 2506 15 2523 23
rect 2506 -23 2523 -15
<< viali >>
rect -2523 -15 -2506 15
rect 2506 -15 2523 15
<< metal1 >>
rect -2526 15 -2503 21
rect -2526 -15 -2523 15
rect -2506 -15 -2503 15
rect -2526 -21 -2503 -15
rect 2503 15 2526 21
rect 2503 -15 2506 15
rect 2523 -15 2526 15
rect 2503 -21 2526 -15
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 50 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_N7YW8T parameters
<< end >>
