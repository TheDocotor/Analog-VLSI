magic
tech sky130A
magscale 1 2
timestamp 1732920865
<< nwell >>
rect -100 -3740 2700 -1600
<< pwell >>
rect -3200 -1600 20200 2400
rect -3200 -3740 -100 -1600
rect 2700 -3740 20200 -1600
rect -3200 -5000 20200 -3740
<< psubdiff >>
rect -3100 2000 -2700 2100
rect -3100 -4600 -3000 2000
rect -2800 -4600 -2700 2000
rect -2600 2000 -2500 2200
rect 19300 2000 19500 2200
rect -2600 1900 19500 2000
rect 19700 1900 20100 2000
rect 19700 -4300 19800 1900
rect 20000 -4300 20100 1900
rect 19700 -4400 20100 -4300
rect -3100 -4700 -2700 -4600
rect -2400 -4600 19600 -4500
rect -2400 -4800 -2300 -4600
rect 19500 -4800 19600 -4600
rect -2400 -4900 19600 -4800
<< nsubdiff >>
rect -40 -1720 1440 -1640
rect 2380 -1720 2640 -1640
rect -40 -3620 60 -1720
rect 2560 -3620 2640 -1720
rect -40 -3700 2660 -3620
<< psubdiffcont >>
rect -3000 -4600 -2800 2000
rect -2500 2000 19300 2200
rect 19800 -4300 20000 1900
rect -2300 -4800 19500 -4600
<< nsubdiffcont >>
rect 1440 -1720 2380 -1640
<< poly >>
rect 9480 -1860 9500 -1780
<< locali >>
rect -3200 2200 20200 2400
rect -3200 2000 -2500 2200
rect 19300 2000 20200 2200
rect -3200 -4600 -3000 2000
rect -2800 1900 20200 2000
rect -2800 1800 19800 1900
rect -2800 -1200 -2600 1800
rect 9600 -20 11560 0
rect 5020 -50 6960 -40
rect 5020 -90 5040 -50
rect 6940 -90 6960 -50
rect 5020 -260 6960 -90
rect 9600 -80 9640 -20
rect 11530 -80 11560 -20
rect 7300 -140 9260 -130
rect 7300 -180 7330 -140
rect 9190 -180 9260 -140
rect 7300 -270 9260 -180
rect 9600 -270 11560 -80
rect -1600 -1085 -1440 -1060
rect -1600 -1200 -1584 -1085
rect -2800 -1482 -1584 -1200
rect -1478 -1200 -1440 -1085
rect -1320 -1085 -1140 -1060
rect -1320 -1200 -1284 -1085
rect -1478 -1482 -1284 -1200
rect -1178 -1200 -1140 -1085
rect -1178 -1482 -400 -1200
rect -2800 -2400 -400 -1482
rect 4820 -1516 4880 -1100
rect 9400 -1270 9460 -1100
rect 9398 -1294 9460 -1270
rect 4820 -1540 5060 -1516
rect 9398 -1520 9458 -1294
rect 4820 -1576 6980 -1540
rect 5000 -1600 6980 -1576
rect 7378 -1580 9458 -1520
rect 7378 -1600 9258 -1580
rect -40 -1720 1440 -1640
rect 2380 -1720 2640 -1640
rect -2800 -4400 -2600 -2400
rect -40 -3620 60 -1720
rect 1218 -3502 1340 -1899
rect 1200 -3510 1340 -3502
rect 1160 -3520 1340 -3510
rect 1160 -3523 1280 -3520
rect 1152 -3552 1280 -3523
rect 1141 -3562 1280 -3552
rect 1141 -3564 1259 -3562
rect 2560 -3620 2640 -1720
rect 7110 -2892 7190 -2440
rect 6140 -2928 8102 -2892
rect 15820 -2940 15880 -1000
rect 19280 -2860 19360 -2300
rect 19280 -2940 19540 -2860
rect -40 -3700 2660 -3620
rect 3370 -3860 3440 -3850
rect 3360 -3890 3440 -3860
rect 3400 -3920 3440 -3890
rect 160 -4400 1130 -4330
rect 1390 -4400 3360 -4320
rect 8260 -4400 8400 -3160
rect 16940 -4400 17100 -3200
rect 19500 -3340 19540 -2940
rect 19600 -4300 19800 1800
rect 20000 -4300 20200 1900
rect 19600 -4400 20200 -4300
rect -2800 -4600 20200 -4400
rect -3200 -4800 -2300 -4600
rect 19500 -4800 20200 -4600
rect -3200 -5000 20200 -4800
<< viali >>
rect -2500 2000 19300 2200
rect -3000 -4600 -2800 2000
rect -1584 293 -1478 690
rect -1284 293 -1178 690
rect 18420 460 18540 520
rect 2318 16 2715 122
rect 4097 16 4494 122
rect 5618 16 6015 122
rect 7397 15 7794 122
rect 12959 114 13356 220
rect 15294 117 15691 223
rect 16019 124 16416 230
rect 18354 127 18751 233
rect -1584 -393 -1478 15
rect -1284 -393 -1178 15
rect 5040 -90 6940 -50
rect 2720 -269 4680 -210
rect 9640 -80 11530 -20
rect 18540 -60 19520 -20
rect 7330 -180 9190 -140
rect 13720 -169 15680 -135
rect 16020 -169 17980 -135
rect -884 -793 -776 -393
rect -584 -793 -476 -393
rect -1584 -1482 -1478 -1085
rect -1284 -1482 -1178 -1085
rect 2540 -1160 2580 -320
rect 2520 -1240 2580 -1160
rect 2540 -1300 2580 -1240
rect 7120 -1300 7160 -320
rect 11700 -1200 11740 -320
rect 13540 -1200 13580 -220
rect 11700 -1260 11750 -1200
rect 11700 -1300 11740 -1260
rect 1440 -1720 2380 -1640
rect 176 -1894 1152 -1860
rect 1412 -1894 2388 -1860
rect 176 -3552 1152 -3518
rect 1412 -3552 2388 -3518
rect 4840 -2640 4880 -1660
rect 9420 -1780 9460 -1660
rect 9420 -1860 9480 -1780
rect 9420 -2640 9460 -1860
rect 18120 -1200 18160 -220
rect 18880 -2340 19200 -2300
rect 160 -3890 1136 -3856
rect 1378 -3890 3354 -3856
rect -260 -4260 -130 -4150
rect 76 -4286 110 -3918
rect 5960 -3960 6000 -2980
rect 14640 -4000 14680 -3020
rect 17400 -3065 19360 -3031
rect 17220 -4100 17260 -3120
rect 19500 -3720 19540 -3480
rect 19800 -4300 20000 1900
rect -2300 -4800 19500 -4600
<< metal1 >>
rect -3200 2200 20200 2400
rect -3200 2000 -2500 2200
rect 19300 2000 20200 2200
rect -3200 -4600 -3000 2000
rect -2800 1900 20200 2000
rect -2800 1800 19800 1900
rect -2800 -1200 -2600 1800
rect -2200 690 18770 1600
rect -2200 400 -1584 690
rect -1620 293 -1584 400
rect -1478 400 -1284 690
rect -1478 293 -1460 400
rect -1620 260 -1460 293
rect -1320 293 -1284 400
rect -1178 520 18770 690
rect -1178 460 18420 520
rect 18540 460 18770 520
rect -1178 400 18770 460
rect -1178 293 -1140 400
rect -1320 280 -1140 293
rect -920 260 -740 400
rect -640 240 -400 400
rect -1620 15 -1440 20
rect -1620 -393 -1584 15
rect -1478 -393 -1440 15
rect -1620 -400 -1440 -393
rect -1340 15 -1120 40
rect -1340 -393 -1284 15
rect -1178 -393 -1120 15
rect -1340 -440 -1120 -393
rect -900 -393 -760 -378
rect -900 -793 -884 -393
rect -776 -793 -760 -393
rect -900 -808 -760 -793
rect -600 -393 -460 -378
rect -600 -793 -584 -393
rect -476 -793 -460 -393
rect -600 -808 -460 -793
rect -1600 -1085 -1440 -1060
rect -1600 -1200 -1584 -1085
rect -2800 -1482 -1584 -1200
rect -1478 -1200 -1440 -1085
rect -1320 -1085 -1140 -1060
rect -1320 -1200 -1284 -1085
rect -1478 -1482 -1284 -1200
rect -1178 -1200 -1140 -1085
rect -1178 -1482 -400 -1200
rect -2800 -2400 -400 -1482
rect 600 -1500 1000 400
rect 2200 172 2600 400
rect 2196 122 2738 172
rect 5600 138 6000 400
rect 12930 238 13370 400
rect 18340 248 18770 400
rect 12930 220 13372 238
rect 2196 16 2318 122
rect 2715 16 2738 122
rect 2196 -18 2738 16
rect 4080 122 4512 138
rect 4080 16 4097 122
rect 4494 16 4512 122
rect 4080 0 4512 16
rect 5600 122 6032 138
rect 5600 16 5618 122
rect 6015 16 6032 122
rect 5600 0 6032 16
rect 7376 122 7942 140
rect 7376 15 7397 122
rect 7794 15 7942 122
rect 12930 114 12959 220
rect 13356 114 13372 220
rect 12930 100 13372 114
rect 15274 223 15706 238
rect 15274 117 15294 223
rect 15691 117 15706 223
rect 15274 100 15706 117
rect 16000 230 16432 248
rect 16000 124 16019 230
rect 16416 124 16432 230
rect 16000 110 16432 124
rect 18334 233 18770 248
rect 18334 127 18354 233
rect 18751 127 18770 233
rect 18334 110 18770 127
rect 7376 2 7942 15
rect 7380 0 7942 2
rect 5600 -2 6030 0
rect 7400 -20 13300 0
rect 7400 -40 9640 -20
rect 4980 -50 9640 -40
rect 4980 -90 5040 -50
rect 6940 -80 9640 -50
rect 11530 -80 13300 -20
rect 6940 -90 13300 -80
rect 4980 -100 13300 -90
rect 7310 -190 7330 -130
rect 9190 -190 9210 -130
rect 2700 -210 4700 -190
rect 2700 -230 2720 -210
rect 2710 -240 2720 -230
rect 4680 -230 4700 -210
rect 13100 -220 13600 -100
rect 15300 -135 15680 100
rect 16000 40 16410 110
rect 16000 -20 19500 40
rect 16000 -60 18540 -20
rect 16000 -130 16410 -60
rect 16000 -135 16412 -130
rect 16000 -168 16020 -135
rect 4680 -240 4690 -230
rect 2480 -1160 2540 -1140
rect 7110 -630 7120 -620
rect 7160 -630 7180 -620
rect 7170 -760 7180 -630
rect 7110 -770 7120 -760
rect 2580 -1150 2600 -1140
rect 2580 -1160 2610 -1150
rect 2480 -1240 2500 -1160
rect 2600 -1240 2610 -1160
rect 2490 -1250 2540 -1240
rect 2580 -1250 2610 -1240
rect 7160 -770 7180 -760
rect 11680 -1190 11700 -1180
rect 11740 -1190 11770 -1180
rect 11680 -1270 11690 -1190
rect 11760 -1270 11770 -1190
rect 13100 -1200 13540 -220
rect 13580 -1200 13600 -220
rect 18110 -220 18180 -200
rect 18110 -1200 18120 -220
rect 18110 -1210 18180 -1200
rect 11680 -1280 11700 -1270
rect 11740 -1280 11770 -1270
rect 600 -1640 2410 -1500
rect -40 -1720 1440 -1640
rect 2380 -1720 2640 -1640
rect -2800 -4400 -2600 -2400
rect -40 -3620 60 -1720
rect 600 -1860 1000 -1720
rect 1410 -1860 2410 -1720
rect 1410 -1894 1412 -1860
rect 2388 -1894 2410 -1860
rect 600 -1900 1000 -1894
rect 1410 -1900 2410 -1894
rect 140 -3500 1160 -3480
rect 140 -3580 160 -3500
rect 140 -3590 1160 -3580
rect 1390 -3510 2410 -3500
rect 1390 -3590 1400 -3510
rect 2400 -3590 2410 -3510
rect 2560 -3620 2640 -1720
rect 4820 -2320 4840 -2120
rect 9470 -1780 9500 -1770
rect 9480 -1860 9500 -1780
rect 4880 -2140 4900 -2120
rect 4880 -2320 4900 -2300
rect 9470 -1880 9500 -1860
rect 18730 -2300 19330 -2290
rect 18730 -2330 18880 -2300
rect 18860 -2340 18880 -2330
rect 19200 -2330 19360 -2300
rect 19200 -2340 19220 -2330
rect 18860 -2360 19220 -2340
rect 19280 -2860 19360 -2330
rect 19280 -2940 19540 -2860
rect 5920 -3000 5960 -2980
rect -40 -3700 2660 -3620
rect 150 -3830 1140 -3820
rect 150 -3890 160 -3830
rect 1360 -3830 3370 -3820
rect 1140 -3890 1150 -3840
rect 1360 -3890 1370 -3830
rect 3360 -3890 3370 -3830
rect 1360 -3900 3370 -3890
rect -320 -4150 76 -3920
rect -320 -4260 -260 -4150
rect -130 -4260 76 -4150
rect -320 -4286 76 -4260
rect 5920 -3960 5940 -3000
rect 6000 -3960 6020 -2980
rect 18390 -3000 18620 -2990
rect 5920 -3980 6020 -3960
rect 14600 -3020 14740 -3000
rect 5960 -4060 6000 -3980
rect 14600 -4000 14620 -3020
rect 14680 -4000 14740 -3020
rect 18390 -3031 18400 -3000
rect 18610 -3031 18620 -3000
rect 18390 -3070 18620 -3065
rect 14600 -4060 14740 -4000
rect 17180 -3960 17220 -3940
rect 19500 -3310 19540 -2940
rect 19490 -3340 19540 -3310
rect 19490 -3460 19530 -3340
rect 19490 -3480 19560 -3460
rect 19490 -3720 19500 -3480
rect 19540 -3720 19560 -3480
rect 19490 -3740 19560 -3720
rect 19490 -3910 19530 -3740
rect 17180 -4080 17200 -3960
rect 17180 -4100 17220 -4080
rect 17260 -4100 17280 -3940
rect -320 -4300 110 -4286
rect 19600 -4300 19800 1800
rect 20000 -4300 20200 1900
rect 19600 -4400 20200 -4300
rect -2800 -4600 20200 -4400
rect -3200 -4800 -2300 -4600
rect 19500 -4800 20200 -4600
rect -3200 -5000 20200 -4800
<< via1 >>
rect 18420 460 18540 520
rect -1584 -393 -1478 15
rect -1284 -393 -1178 15
rect -884 -793 -776 -393
rect -584 -793 -476 -393
rect 4097 16 4494 122
rect 7330 -140 9190 -130
rect 7330 -180 9190 -140
rect 7330 -190 9190 -180
rect 2720 -269 4680 -210
rect 7110 -760 7120 -630
rect 7120 -760 7160 -630
rect 7160 -760 7170 -630
rect 2500 -1240 2520 -1160
rect 2520 -1240 2580 -1160
rect 2580 -1240 2600 -1160
rect 11690 -1270 11700 -1190
rect 11700 -1200 11740 -1190
rect 11740 -1200 11760 -1190
rect 11700 -1260 11750 -1200
rect 11750 -1260 11760 -1200
rect 11700 -1270 11740 -1260
rect 11740 -1270 11760 -1260
rect 18120 -1200 18160 -220
rect 18160 -1200 18180 -220
rect 160 -3518 1160 -3500
rect 160 -3552 176 -3518
rect 176 -3552 1152 -3518
rect 1152 -3552 1160 -3518
rect 160 -3580 1160 -3552
rect 1400 -3518 2400 -3510
rect 1400 -3552 1412 -3518
rect 1412 -3552 2388 -3518
rect 2388 -3552 2400 -3518
rect 1400 -3590 2400 -3552
rect 9420 -1860 9480 -1780
rect 4840 -2300 4880 -2140
rect 4880 -2300 4900 -2140
rect 160 -3856 1140 -3830
rect 160 -3890 1136 -3856
rect 1136 -3890 1140 -3856
rect 1370 -3856 3360 -3830
rect 1370 -3890 1378 -3856
rect 1378 -3890 3354 -3856
rect 3354 -3890 3360 -3856
rect -260 -4260 -130 -4150
rect 5940 -3960 5960 -3000
rect 5960 -3960 6000 -3000
rect 14620 -4000 14640 -3020
rect 14640 -4000 14680 -3020
rect 18400 -3031 18610 -3000
rect 18400 -3060 18610 -3031
rect 17200 -4080 17220 -3960
rect 17220 -4080 17260 -3960
<< metal2 >>
rect -1600 500 1300 700
rect -1600 30 -1400 500
rect -1620 15 -1400 30
rect -1620 -393 -1584 15
rect -1478 0 -1400 15
rect -1340 15 -1120 40
rect -1478 -393 -1440 0
rect -1620 -410 -1440 -393
rect -1340 -393 -1284 15
rect -1178 0 -1120 15
rect -1178 -200 500 0
rect -1178 -393 -1120 -200
rect -1340 -440 -1120 -393
rect -932 -393 -706 -366
rect -932 -793 -884 -393
rect -776 -793 -706 -393
rect -932 -2140 -706 -793
rect -620 -393 -440 -360
rect -620 -793 -584 -393
rect -476 -793 -440 -393
rect -620 -1780 -440 -793
rect 300 -1100 500 -200
rect 1100 -600 1300 500
rect 18380 520 18620 560
rect 18380 460 18420 520
rect 18540 460 18620 520
rect 4080 140 4520 160
rect 4080 122 4530 140
rect 4080 16 4097 122
rect 4494 16 4530 122
rect 4080 -70 4530 16
rect 4080 -100 9260 -70
rect 4080 -130 18240 -100
rect 4080 -170 7330 -130
rect 4080 -200 4530 -170
rect 7310 -190 7330 -170
rect 9190 -190 18240 -130
rect 7310 -200 18240 -190
rect 2710 -210 4690 -200
rect 2710 -269 2720 -210
rect 4680 -269 4690 -210
rect 2710 -270 4690 -269
rect 18110 -220 18240 -200
rect 1100 -630 7200 -600
rect 1100 -760 7110 -630
rect 7170 -760 7200 -630
rect 1100 -800 7200 -760
rect 300 -1160 11800 -1100
rect 300 -1240 2500 -1160
rect 2600 -1190 11800 -1160
rect 2600 -1240 11690 -1190
rect 300 -1270 11690 -1240
rect 11760 -1270 11800 -1190
rect 18110 -1200 18120 -220
rect 18180 -1200 18240 -220
rect 18110 -1210 18240 -1200
rect 300 -1300 11800 -1270
rect -620 -1860 9420 -1780
rect 9480 -1860 9490 -1780
rect -620 -2020 -440 -1860
rect 9410 -1880 9490 -1860
rect 4820 -2140 4920 -2120
rect -952 -2300 4840 -2140
rect 4900 -2300 4920 -2140
rect -952 -2302 4920 -2300
rect 4820 -2320 4920 -2302
rect 18380 -3000 18620 460
rect 140 -3500 1180 -3480
rect 140 -3580 160 -3500
rect 1160 -3580 1180 -3500
rect 140 -3600 1180 -3580
rect 1380 -3510 2430 -3490
rect 1380 -3590 1400 -3510
rect 2400 -3590 2430 -3510
rect 1380 -3600 2430 -3590
rect 170 -3820 1080 -3600
rect 1410 -3820 2430 -3600
rect 3020 -3820 5940 -3000
rect 140 -3830 1150 -3820
rect 140 -3890 160 -3830
rect 1140 -3890 1150 -3830
rect 140 -3900 1150 -3890
rect 1360 -3830 5940 -3820
rect 1360 -3890 1370 -3830
rect 3360 -3890 5940 -3830
rect 1360 -3900 3370 -3890
rect 3660 -3960 5940 -3890
rect 6000 -3002 14640 -3000
rect 6000 -3020 14696 -3002
rect 6000 -3960 14620 -3020
rect 3660 -4000 14620 -3960
rect 14680 -4000 14696 -3020
rect 18380 -3060 18400 -3000
rect 18610 -3060 18620 -3000
rect 18380 -3080 18620 -3060
rect 3660 -4060 14696 -4000
rect 17180 -3960 17280 -3940
rect 17180 -4080 17200 -3960
rect 17260 -4080 17280 -3960
rect 17180 -4100 17280 -4080
rect -280 -4150 -80 -4120
rect -280 -4260 -260 -4150
rect -130 -4200 -80 -4150
rect 17200 -4200 17260 -4100
rect -130 -4260 17260 -4200
rect -280 -4280 17260 -4260
rect -200 -4400 17260 -4280
use Gilbert  Gilbert_0
timestamp 1732917019
transform 0 1 4800 -1 0 -100
box 0 -2300 1404 2400
use Gilbert  Gilbert_1
timestamp 1732917019
transform 0 1 9380 -1 0 -100
box 0 -2300 1404 2400
use Gilbert  Gilbert_2
timestamp 1732917019
transform 0 1 7100 -1 0 -1440
box 0 -2300 1404 2400
use Gilbert  Gilbert_3
timestamp 1732917019
transform 0 1 15800 -1 0 0
box 0 -2300 1404 2400
use if_res  if_res_0
timestamp 1729706060
transform 0 1 12940 -1 0 -162
box -400 0 -262 2766
use if_res  if_res_1
timestamp 1729706060
transform 0 1 16000 -1 0 -152
box -400 0 -262 2766
use LOp_resistor  LOp_resistor_0
timestamp 1729706114
transform 1 0 -1400 0 1 -1000
box -200 -500 -52 1708
use LOp_resistor  LOp_resistor_1
timestamp 1729706114
transform 1 0 -1100 0 1 -1000
box -200 -500 -52 1708
use nmos_40  nmos_40_0
timestamp 1732917019
transform 0 -1 8520 -1 0 -4160
box -1400 200 0 2600
use nmos_40  nmos_40_1
timestamp 1732917019
transform 0 -1 19780 1 0 -2920
box -1400 200 0 2600
use nmos_40  nmos_40_2
timestamp 1732917019
transform 0 -1 17200 -1 0 -4200
box -1400 200 0 2600
use nmos_40  nmos_40_3
timestamp 1732917019
transform -1 0 18340 0 1 -2580
box -1400 200 0 2600
use sky130_fd_pr__nfet_01v8_8WUFR5  sky130_fd_pr__nfet_01v8_8WUFR5_0
timestamp 1732920865
transform 0 -1 617 -1 0 -4102
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_P82RFK  sky130_fd_pr__nfet_01v8_P82RFK_0
timestamp 1732920865
transform 0 1 2397 -1 0 -4102
box -258 -1057 258 1057
use sky130_fd_pr__pfet_01v8_AXDRNP  sky130_fd_pr__pfet_01v8_AXDRNP_0
timestamp 1732122809
transform 0 -1 1864 -1 0 -2706
box -894 -598 894 564
use sky130_fd_pr__pfet_01v8_GXDZBM  sky130_fd_pr__pfet_01v8_GXDZBM_1
timestamp 1732122809
transform 0 1 700 -1 0 -2706
box -894 -598 894 564
use Vdd_res  Vdd_res_0
timestamp 1729706186
transform 0 1 2300 -1 0 138
box 0 0 138 2212
use Vdd_res  Vdd_res_1
timestamp 1729706186
transform 0 1 5600 -1 0 138
box 0 0 138 2212
<< labels >>
flabel metal1 -700 -4900 -700 -4900 0 FreeSans 1600 0 0 0 VSS
port 8 nsew
flabel metal1 -1200 -100 -1200 -100 0 FreeSans 1600 0 0 0 LOp
port 2 nsew
flabel via1 -500 -600 -500 -600 0 FreeSans 1600 0 0 0 RFn
port 5 nsew
flabel via1 -800 -700 -800 -700 0 FreeSans 1600 0 0 0 RFp
port 4 nsew
flabel viali 7608 82 7610 84 0 FreeSans 1600 0 0 0 IF--
flabel via1 4328 70 4328 70 0 FreeSans 1600 0 0 0 IF++
flabel metal1 3000 1100 3000 1100 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel locali 15848 -2038 15848 -2038 0 FreeSans 1600 0 0 0 Vamp
flabel locali 7144 -2614 7144 -2614 0 FreeSans 1600 0 0 0 Vbottom
flabel locali 9432 -1360 9432 -1360 0 FreeSans 1600 0 0 0 Vmid2
flabel locali 4852 -1364 4852 -1364 0 FreeSans 1600 0 0 0 Vmid
flabel metal1 -1520 -240 -1520 -240 0 FreeSans 1600 0 0 0 LOn
port 3 nsew
flabel metal1 -140 -4100 -140 -4100 0 FreeSans 1600 0 0 0 Vref
port 7 nsew
flabel viali 15480 160 15480 160 0 FreeSans 1600 0 0 0 IFp
flabel viali 16200 180 16200 180 0 FreeSans 1600 0 0 0 IFn
flabel metal1 19320 -2580 19320 -2580 0 FreeSans 1600 0 0 0 IF
port 1 nsew
flabel via1 5980 -3520 5980 -3520 0 FreeSans 1600 0 0 0 VM
port 6 nsew
<< end >>
