magic
tech sky130A
timestamp 1728490836
<< pwell >>
rect -341 -605 341 605
<< nmos >>
rect -243 -500 -143 500
rect -114 -500 -14 500
rect 14 -500 114 500
rect 143 -500 243 500
<< ndiff >>
rect -272 494 -243 500
rect -272 -494 -266 494
rect -249 -494 -243 494
rect -272 -500 -243 -494
rect -143 494 -114 500
rect -143 -494 -137 494
rect -120 -494 -114 494
rect -143 -500 -114 -494
rect -14 494 14 500
rect -14 -494 -8 494
rect 8 -494 14 494
rect -14 -500 14 -494
rect 114 494 143 500
rect 114 -494 120 494
rect 137 -494 143 494
rect 114 -500 143 -494
rect 243 494 272 500
rect 243 -494 249 494
rect 266 -494 272 494
rect 243 -500 272 -494
<< ndiffc >>
rect -266 -494 -249 494
rect -137 -494 -120 494
rect -8 -494 8 494
rect 120 -494 137 494
rect 249 -494 266 494
<< psubdiff >>
rect -323 570 -275 587
rect 275 570 323 587
rect -323 539 -306 570
rect 306 539 323 570
rect -323 -570 -306 -539
rect 306 -570 323 -539
rect -323 -587 -275 -570
rect 275 -587 323 -570
<< psubdiffcont >>
rect -275 570 275 587
rect -323 -539 -306 539
rect 306 -539 323 539
rect -275 -587 275 -570
<< poly >>
rect -243 536 -143 544
rect -243 519 -235 536
rect -151 519 -143 536
rect -243 500 -143 519
rect -114 536 -14 544
rect -114 519 -106 536
rect -22 519 -14 536
rect -114 500 -14 519
rect 14 536 114 544
rect 14 519 22 536
rect 106 519 114 536
rect 14 500 114 519
rect 143 536 243 544
rect 143 519 151 536
rect 235 519 243 536
rect 143 500 243 519
rect -243 -519 -143 -500
rect -243 -536 -235 -519
rect -151 -536 -143 -519
rect -243 -544 -143 -536
rect -114 -519 -14 -500
rect -114 -536 -106 -519
rect -22 -536 -14 -519
rect -114 -544 -14 -536
rect 14 -519 114 -500
rect 14 -536 22 -519
rect 106 -536 114 -519
rect 14 -544 114 -536
rect 143 -519 243 -500
rect 143 -536 151 -519
rect 235 -536 243 -519
rect 143 -544 243 -536
<< polycont >>
rect -235 519 -151 536
rect -106 519 -22 536
rect 22 519 106 536
rect 151 519 235 536
rect -235 -536 -151 -519
rect -106 -536 -22 -519
rect 22 -536 106 -519
rect 151 -536 235 -519
<< locali >>
rect -323 570 -275 587
rect 275 570 323 587
rect -323 539 -306 570
rect 306 539 323 570
rect -243 519 -235 536
rect -151 519 -143 536
rect -114 519 -106 536
rect -22 519 -14 536
rect 14 519 22 536
rect 106 519 114 536
rect 143 519 151 536
rect 235 519 243 536
rect -266 494 -249 502
rect -266 -502 -249 -494
rect -137 494 -120 502
rect -137 -502 -120 -494
rect -8 494 8 502
rect -8 -502 8 -494
rect 120 494 137 502
rect 120 -502 137 -494
rect 249 494 266 502
rect 249 -502 266 -494
rect -243 -536 -235 -519
rect -151 -536 -143 -519
rect -114 -536 -106 -519
rect -22 -536 -14 -519
rect 14 -536 22 -519
rect 106 -536 114 -519
rect 143 -536 151 -519
rect 235 -536 243 -519
rect -323 -570 -306 -539
rect 306 -570 323 -539
rect -323 -587 -275 -570
rect 275 -587 323 -570
<< viali >>
rect -235 519 -151 536
rect -106 519 -22 536
rect 22 519 106 536
rect 151 519 235 536
rect -266 -494 -249 494
rect -137 -494 -120 494
rect -8 -494 8 494
rect 120 -494 137 494
rect 249 -494 266 494
rect -235 -536 -151 -519
rect -106 -536 -22 -519
rect 22 -536 106 -519
rect 151 -536 235 -519
<< metal1 >>
rect -241 536 -145 539
rect -241 519 -235 536
rect -151 519 -145 536
rect -241 516 -145 519
rect -112 536 -16 539
rect -112 519 -106 536
rect -22 519 -16 536
rect -112 516 -16 519
rect 16 536 112 539
rect 16 519 22 536
rect 106 519 112 536
rect 16 516 112 519
rect 145 536 241 539
rect 145 519 151 536
rect 235 519 241 536
rect 145 516 241 519
rect -269 494 -246 500
rect -269 -494 -266 494
rect -249 -494 -246 494
rect -269 -500 -246 -494
rect -140 494 -117 500
rect -140 -494 -137 494
rect -120 -494 -117 494
rect -140 -500 -117 -494
rect -11 494 11 500
rect -11 -494 -8 494
rect 8 -494 11 494
rect -11 -500 11 -494
rect 117 494 140 500
rect 117 -494 120 494
rect 137 -494 140 494
rect 117 -500 140 -494
rect 246 494 269 500
rect 246 -494 249 494
rect 266 -494 269 494
rect 246 -500 269 -494
rect -241 -519 -145 -516
rect -241 -536 -235 -519
rect -151 -536 -145 -519
rect -241 -539 -145 -536
rect -112 -519 -16 -516
rect -112 -536 -106 -519
rect -22 -536 -16 -519
rect -112 -539 -16 -536
rect 16 -519 112 -516
rect 16 -536 22 -519
rect 106 -536 112 -519
rect 16 -539 112 -536
rect 145 -519 241 -516
rect 145 -536 151 -519
rect 235 -536 241 -519
rect 145 -539 241 -536
<< properties >>
string FIXED_BBOX -315 -578 315 578
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_TCXCTP parameters
<< end >>
