magic
tech sky130A
timestamp 1729287489
<< pwell >>
rect -348 -155 348 155
<< nmos >>
rect -250 -50 250 50
<< ndiff >>
rect -279 44 -250 50
rect -279 -44 -273 44
rect -256 -44 -250 44
rect -279 -50 -250 -44
rect 250 44 279 50
rect 250 -44 256 44
rect 273 -44 279 44
rect 250 -50 279 -44
<< ndiffc >>
rect -273 -44 -256 44
rect 256 -44 273 44
<< psubdiff >>
rect -330 120 -282 137
rect 282 120 330 137
rect -330 89 -313 120
rect 313 89 330 120
rect -330 -120 -313 -89
rect 313 -120 330 -89
rect -330 -137 -282 -120
rect 282 -137 330 -120
<< psubdiffcont >>
rect -282 120 282 137
rect -330 -89 -313 89
rect 313 -89 330 89
rect -282 -137 282 -120
<< poly >>
rect -250 86 250 94
rect -250 69 -242 86
rect 242 69 250 86
rect -250 50 250 69
rect -250 -69 250 -50
rect -250 -86 -242 -69
rect 242 -86 250 -69
rect -250 -94 250 -86
<< polycont >>
rect -242 69 242 86
rect -242 -86 242 -69
<< locali >>
rect -330 120 -282 137
rect 282 120 330 137
rect -330 89 -313 120
rect 313 89 330 120
rect -250 69 -242 86
rect 242 69 250 86
rect -273 44 -256 52
rect -273 -52 -256 -44
rect 256 44 273 52
rect 256 -52 273 -44
rect -250 -86 -242 -69
rect 242 -86 250 -69
rect -330 -120 -313 -89
rect 313 -120 330 -89
rect -330 -137 -282 -120
rect 282 -137 330 -120
<< viali >>
rect -242 69 242 86
rect -273 -44 -256 44
rect 256 -44 273 44
rect -242 -86 242 -69
<< metal1 >>
rect -248 86 248 89
rect -248 69 -242 86
rect 242 69 248 86
rect -248 66 248 69
rect -276 44 -253 50
rect -276 -44 -273 44
rect -256 -44 -253 44
rect -276 -50 -253 -44
rect 253 44 276 50
rect 253 -44 256 44
rect 273 -44 276 44
rect 253 -50 276 -44
rect -248 -69 248 -66
rect -248 -86 -242 -69
rect 242 -86 248 -69
rect -248 -89 248 -86
<< properties >>
string FIXED_BBOX -321 -128 321 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_4HNDKD parameters
<< end >>
