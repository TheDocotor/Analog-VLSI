** sch_path: /home/renslow/Documents/ece5120/hw02/xschem/cs_amp.sch
**.subckt cs_amp VDD Vo Vin VSS
*.ipin Vin
*.ipin VDD
*.opin Vo
*.ipin VSS
x1 V_D V_gate net1 VSS my_nmos
C1 Vin V_gate 100u m=1
C2 Vo V_D 100u m=1
Vmeas net1 VSS 0
.save i(vmeas)
R1 VDD V_gate 10k m=1
R2 V_gate VSS 12.5k m=1
R3 VDD V_D 3.73k m=1
**.ends
.end
