magic
tech sky130A
timestamp 1731517815
<< pwell >>
rect -1325 -950 0 250
<< nmos >>
rect -1000 0 -200 100
rect -1000 -200 -200 -100
rect -1000 -400 -200 -300
rect -1000 -600 -200 -500
rect -1000 -800 -200 -700
<< ndiff >>
rect -1000 175 -200 200
rect -1000 125 -975 175
rect -225 125 -200 175
rect -1000 100 -200 125
rect -1000 -25 -200 0
rect -1000 -75 -975 -25
rect -225 -75 -200 -25
rect -1000 -100 -200 -75
rect -1000 -225 -200 -200
rect -1000 -275 -975 -225
rect -225 -275 -200 -225
rect -1000 -300 -200 -275
rect -1000 -425 -200 -400
rect -1000 -475 -975 -425
rect -225 -475 -200 -425
rect -1000 -500 -200 -475
rect -1000 -625 -200 -600
rect -1000 -675 -975 -625
rect -225 -675 -200 -625
rect -1000 -700 -200 -675
rect -1000 -825 -200 -800
rect -1000 -875 -975 -825
rect -225 -875 -200 -825
rect -1000 -900 -200 -875
<< ndiffc >>
rect -975 125 -225 175
rect -975 -75 -225 -25
rect -975 -275 -225 -225
rect -975 -475 -225 -425
rect -975 -675 -225 -625
rect -975 -875 -225 -825
<< poly >>
rect -1300 75 -1000 100
rect -1300 -775 -1275 75
rect -1225 0 -1000 75
rect -200 0 -100 100
rect -1225 -100 -1100 0
rect -1225 -200 -1000 -100
rect -200 -200 -100 -100
rect -1225 -300 -1100 -200
rect -1225 -400 -1000 -300
rect -200 -400 -100 -300
rect -1225 -500 -1100 -400
rect -1225 -600 -1000 -500
rect -200 -600 -100 -500
rect -1225 -700 -1100 -600
rect -1225 -775 -1000 -700
rect -1300 -800 -1000 -775
rect -200 -800 -100 -700
<< polycont >>
rect -1275 -775 -1225 75
<< locali >>
rect -1000 175 -25 200
rect -1000 125 -975 175
rect -225 125 -25 175
rect -1000 100 -25 125
rect -1300 75 -1200 100
rect -1300 -775 -1275 75
rect -1225 -775 -1200 75
rect -1300 -800 -1200 -775
rect -1150 -25 -200 0
rect -1150 -75 -975 -25
rect -225 -75 -200 -25
rect -1150 -100 -200 -75
rect -1150 -400 -1050 -100
rect -125 -200 -25 100
rect -1000 -225 -25 -200
rect -1000 -275 -975 -225
rect -225 -275 -25 -225
rect -1000 -300 -25 -275
rect -1150 -425 -200 -400
rect -1150 -475 -975 -425
rect -225 -475 -200 -425
rect -1150 -500 -200 -475
rect -1150 -800 -1050 -500
rect -125 -600 -25 -300
rect -1000 -625 -25 -600
rect -1000 -675 -975 -625
rect -225 -675 -25 -625
rect -1000 -700 -25 -675
rect -1150 -825 -200 -800
rect -1150 -875 -975 -825
rect -225 -875 -200 -825
rect -1150 -900 -200 -875
<< labels >>
flabel ndiffc -750 150 -750 150 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel polycont -1250 -300 -1250 -300 0 FreeSans 800 0 0 0 G
port 1 nsew
flabel ndiffc -750 -850 -750 -850 0 FreeSans 800 0 0 0 S
port 2 nsew
flabel pwell -1200 175 -1200 175 0 FreeSans 800 0 0 0 B
port 3 nsew
<< end >>
