magic
tech sky130A
timestamp 1726935614
<< pwell >>
rect -1153 -49 -454 1146
<< nmos >>
rect -1040 52 -565 1038
<< ndiff >>
rect -1076 1007 -1040 1038
rect -1076 84 -1067 1007
rect -1049 84 -1040 1007
rect -1076 52 -1040 84
rect -565 989 -525 1038
rect -565 77 -553 989
rect -536 77 -525 989
rect -565 52 -525 77
<< ndiffc >>
rect -1067 84 -1049 1007
rect -553 77 -536 989
<< psubdiff >>
rect -1133 1101 -1076 1124
rect -521 1101 -473 1124
rect -1133 1070 -1111 1101
rect -490 1065 -473 1101
rect -1133 -13 -1111 15
rect -490 -13 -473 29
rect -1133 -30 -1068 -13
rect -521 -30 -473 -13
<< psubdiffcont >>
rect -1076 1101 -521 1124
rect -1133 15 -1111 1070
rect -490 29 -473 1065
rect -1068 -30 -521 -13
<< poly >>
rect -1040 1074 -565 1083
rect -1040 1057 -1022 1074
rect -577 1057 -565 1074
rect -1040 1038 -565 1057
rect -1040 33 -565 52
rect -1040 16 -1022 33
rect -577 16 -565 33
rect -1040 5 -565 16
<< polycont >>
rect -1022 1057 -577 1074
rect -1022 16 -577 33
<< locali >>
rect -1131 1122 -1076 1124
rect -1133 1101 -1076 1122
rect -521 1101 -473 1124
rect -1133 1070 -1111 1101
rect -1040 1057 -1022 1074
rect -577 1057 -565 1074
rect -490 1065 -473 1101
rect -1067 1007 -1049 1038
rect -1067 49 -1049 84
rect -553 989 -535 1037
rect -536 77 -535 989
rect -553 52 -535 77
rect -1040 16 -1022 33
rect -577 16 -565 33
rect -1133 -13 -1111 15
rect -490 -13 -473 29
rect -1133 -30 -1068 -13
rect -521 -30 -473 -13
<< viali >>
rect -1022 1057 -577 1074
rect -1067 84 -1049 1007
rect -553 77 -536 989
rect -1022 16 -577 33
<< metal1 >>
rect -1036 1074 -570 1078
rect -1036 1057 -1022 1074
rect -577 1057 -570 1074
rect -1036 1050 -570 1057
rect -1071 1007 -1045 1038
rect -1071 84 -1067 1007
rect -1049 84 -1045 1007
rect -1071 52 -1045 84
rect -558 989 -530 1038
rect -558 77 -553 989
rect -536 77 -530 989
rect -558 52 -530 77
rect -1032 33 -570 38
rect -1032 16 -1022 33
rect -577 16 -570 33
rect -1032 13 -570 16
<< labels >>
flabel viali -1056 557 -1056 557 0 FreeSans 200 0 0 0 D
port 0 nsew
flabel viali -812 1066 -812 1066 0 FreeSans 200 0 0 0 G
port 1 nsew
flabel viali -546 562 -546 562 0 FreeSans 200 0 0 0 S
port 2 nsew
flabel psubdiffcont -809 1111 -809 1111 0 FreeSans 200 0 0 0 B
port 3 nsew
<< end >>
