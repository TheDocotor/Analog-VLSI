magic
tech sky130A
timestamp 1731516743
<< pwell >>
rect -900 -1100 900 600
<< nmos >>
rect -400 300 600 400
rect -400 100 600 200
rect -400 -100 600 0
rect -400 -300 600 -200
rect -400 -500 600 -400
rect -400 -700 600 -600
rect -400 -900 600 -800
<< ndiff >>
rect -400 475 600 500
rect -400 425 -375 475
rect 575 425 600 475
rect -400 400 600 425
rect -400 275 600 300
rect -400 225 -375 275
rect 575 225 600 275
rect -400 200 600 225
rect -400 75 600 100
rect -400 25 -375 75
rect 575 25 600 75
rect -400 0 600 25
rect -400 -125 600 -100
rect -400 -175 -375 -125
rect 575 -175 600 -125
rect -400 -200 600 -175
rect -400 -325 600 -300
rect -400 -375 -375 -325
rect 575 -375 600 -325
rect -400 -400 600 -375
rect -400 -525 600 -500
rect -400 -575 -375 -525
rect 575 -575 600 -525
rect -400 -600 600 -575
rect -400 -725 600 -700
rect -400 -775 -375 -725
rect 575 -775 600 -725
rect -400 -800 600 -775
rect -400 -925 600 -900
rect -400 -975 -375 -925
rect 575 -975 600 -925
rect -400 -1000 600 -975
<< ndiffc >>
rect -375 425 575 475
rect -375 225 575 275
rect -375 25 575 75
rect -375 -175 575 -125
rect -375 -375 575 -325
rect -375 -575 575 -525
rect -375 -775 575 -725
rect -375 -975 575 -925
<< poly >>
rect -700 375 -400 400
rect -700 -875 -675 375
rect -625 300 -400 375
rect 600 300 700 400
rect -625 200 -550 300
rect -625 100 -400 200
rect 600 100 700 200
rect -625 0 -550 100
rect -625 -100 -400 0
rect 600 -100 700 0
rect -625 -200 -550 -100
rect -625 -300 -400 -200
rect 600 -300 700 -200
rect -625 -400 -550 -300
rect -625 -500 -400 -400
rect 600 -500 700 -400
rect -625 -600 -550 -500
rect -625 -700 -400 -600
rect 600 -700 700 -600
rect -625 -800 -550 -700
rect -625 -875 -400 -800
rect -700 -900 -400 -875
rect 600 -900 700 -800
<< polycont >>
rect -675 -875 -625 375
<< locali >>
rect -550 475 600 500
rect -550 425 -375 475
rect 575 425 600 475
rect -550 400 600 425
rect -700 375 -600 400
rect -700 -875 -675 375
rect -625 -875 -600 375
rect -550 100 -450 400
rect -400 275 750 300
rect -400 225 -375 275
rect 575 225 750 275
rect -400 200 750 225
rect -550 75 600 100
rect -550 25 -375 75
rect 575 25 600 75
rect -550 0 600 25
rect -550 -300 -450 0
rect 650 -100 750 200
rect -400 -125 750 -100
rect -400 -175 -375 -125
rect 575 -175 750 -125
rect -400 -200 750 -175
rect -550 -325 600 -300
rect -550 -375 -375 -325
rect 575 -375 600 -325
rect -550 -400 600 -375
rect -550 -700 -450 -400
rect 650 -500 750 -200
rect -400 -525 750 -500
rect -400 -575 -375 -525
rect 575 -575 750 -525
rect -400 -600 750 -575
rect -550 -725 600 -700
rect -550 -775 -375 -725
rect 575 -775 600 -725
rect -550 -800 600 -775
rect -700 -900 -600 -875
rect 650 -900 750 -600
rect -400 -925 750 -900
rect -400 -975 -375 -925
rect 575 -975 750 -925
rect -400 -1000 750 -975
<< labels >>
flabel ndiffc 100 450 100 450 0 FreeSans 400 0 0 0 D
port 0 nsew
flabel polycont -650 -275 -650 -275 0 FreeSans 400 0 0 0 G
port 1 nsew
flabel ndiffc 100 -950 100 -950 0 FreeSans 400 0 0 0 S
port 2 nsew
flabel pwell -775 500 -775 500 0 FreeSans 400 0 0 0 B
port 3 nsew
<< end >>
