magic
tech sky130A
magscale 1 2
timestamp 1730311536
<< nwell >>
rect 250 1547 2650 1550
rect 234 -468 2665 1547
<< nsubdiff >>
rect 273 1495 2626 1508
rect 273 -403 299 1495
rect 338 1430 2561 1456
rect 338 -351 351 1430
rect 2548 -351 2561 1430
rect 338 -364 2561 -351
rect 2600 -403 2626 1495
rect 273 -429 2626 -403
<< nsubdiffcont >>
rect 299 1456 2600 1495
rect 299 -364 338 1456
rect 2561 -364 2600 1456
rect 299 -403 2600 -364
<< locali >>
rect 273 1495 2626 1508
rect 273 -403 299 1495
rect 338 1430 2561 1456
rect 338 -351 351 1430
rect 2548 -351 2561 1430
rect 338 -364 2561 -351
rect 2600 -403 2626 1495
rect 273 -429 2626 -403
<< viali >>
rect 750 -225 1300 -175
rect 1600 -225 2150 -175
rect 750 -675 1300 -625
rect 1600 -675 2150 -625
<< metal1 >>
rect 725 -175 1325 -150
rect 725 -225 750 -175
rect 1300 -225 1325 -175
rect 725 -625 1325 -225
rect 725 -675 750 -625
rect 1300 -675 1325 -625
rect 725 -700 1325 -675
rect 1575 -175 2175 -150
rect 1575 -225 1600 -175
rect 2150 -225 2175 -175
rect 1575 -625 2175 -225
rect 1575 -675 1600 -625
rect 2150 -675 2175 -625
rect 1575 -700 2175 -675
use n20x1  n20x1_1
timestamp 1730304573
transform -1 0 2475 0 1 -1100
box -100 -1200 1200 600
use n20x1  n20x1_2
timestamp 1730304573
transform 1 0 425 0 1 -1100
box -100 -1200 1200 600
use p20x1  p20x1_0
timestamp 1730302828
transform 1 0 425 0 -1 250
box -25 -1150 1075 550
use p20x1  p20x1_1
timestamp 1730302828
transform -1 0 2475 0 -1 250
box -25 -1150 1075 550
<< end >>
