magic
tech sky130A
magscale 1 2
timestamp 1728490836
<< pwell >>
rect -683 -1210 683 1210
<< nmos >>
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
<< ndiff >>
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
<< ndiffc >>
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
<< psubdiff >>
rect -647 1140 -551 1174
rect 551 1140 647 1174
rect -647 1078 -613 1140
rect 613 1078 647 1140
rect -647 -1140 -613 -1078
rect 613 -1140 647 -1078
rect -647 -1174 -551 -1140
rect 551 -1174 647 -1140
<< psubdiffcont >>
rect -551 1140 551 1174
rect -647 -1078 -613 1078
rect 613 -1078 647 1078
rect -551 -1174 551 -1140
<< poly >>
rect -487 1072 -287 1088
rect -487 1038 -471 1072
rect -303 1038 -287 1072
rect -487 1000 -287 1038
rect -229 1072 -29 1088
rect -229 1038 -213 1072
rect -45 1038 -29 1072
rect -229 1000 -29 1038
rect 29 1072 229 1088
rect 29 1038 45 1072
rect 213 1038 229 1072
rect 29 1000 229 1038
rect 287 1072 487 1088
rect 287 1038 303 1072
rect 471 1038 487 1072
rect 287 1000 487 1038
rect -487 -1038 -287 -1000
rect -487 -1072 -471 -1038
rect -303 -1072 -287 -1038
rect -487 -1088 -287 -1072
rect -229 -1038 -29 -1000
rect -229 -1072 -213 -1038
rect -45 -1072 -29 -1038
rect -229 -1088 -29 -1072
rect 29 -1038 229 -1000
rect 29 -1072 45 -1038
rect 213 -1072 229 -1038
rect 29 -1088 229 -1072
rect 287 -1038 487 -1000
rect 287 -1072 303 -1038
rect 471 -1072 487 -1038
rect 287 -1088 487 -1072
<< polycont >>
rect -471 1038 -303 1072
rect -213 1038 -45 1072
rect 45 1038 213 1072
rect 303 1038 471 1072
rect -471 -1072 -303 -1038
rect -213 -1072 -45 -1038
rect 45 -1072 213 -1038
rect 303 -1072 471 -1038
<< locali >>
rect -647 1140 -551 1174
rect 551 1140 647 1174
rect -647 1078 -613 1140
rect 613 1078 647 1140
rect -487 1038 -471 1072
rect -303 1038 -287 1072
rect -229 1038 -213 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 213 1038 229 1072
rect 287 1038 303 1072
rect 471 1038 487 1072
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect -487 -1072 -471 -1038
rect -303 -1072 -287 -1038
rect -229 -1072 -213 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 213 -1072 229 -1038
rect 287 -1072 303 -1038
rect 471 -1072 487 -1038
rect -647 -1140 -613 -1078
rect 613 -1140 647 -1078
rect -647 -1174 -551 -1140
rect 551 -1174 647 -1140
<< viali >>
rect -471 1038 -303 1072
rect -213 1038 -45 1072
rect 45 1038 213 1072
rect 303 1038 471 1072
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect -471 -1072 -303 -1038
rect -213 -1072 -45 -1038
rect 45 -1072 213 -1038
rect 303 -1072 471 -1038
<< metal1 >>
rect -483 1072 -291 1078
rect -483 1038 -471 1072
rect -303 1038 -291 1072
rect -483 1032 -291 1038
rect -225 1072 -33 1078
rect -225 1038 -213 1072
rect -45 1038 -33 1072
rect -225 1032 -33 1038
rect 33 1072 225 1078
rect 33 1038 45 1072
rect 213 1038 225 1072
rect 33 1032 225 1038
rect 291 1072 483 1078
rect 291 1038 303 1072
rect 471 1038 483 1072
rect 291 1032 483 1038
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect -483 -1038 -291 -1032
rect -483 -1072 -471 -1038
rect -303 -1072 -291 -1038
rect -483 -1078 -291 -1072
rect -225 -1038 -33 -1032
rect -225 -1072 -213 -1038
rect -45 -1072 -33 -1038
rect -225 -1078 -33 -1072
rect 33 -1038 225 -1032
rect 33 -1072 45 -1038
rect 213 -1072 225 -1038
rect 33 -1078 225 -1072
rect 291 -1038 483 -1032
rect 291 -1072 303 -1038
rect 471 -1072 483 -1038
rect 291 -1078 483 -1072
<< properties >>
string FIXED_BBOX -630 -1157 630 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_01v8_TCXCTP parameters
<< end >>
