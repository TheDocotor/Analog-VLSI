magic
tech sky130A
timestamp 1732735011
<< pwell >>
rect 240 -1020 450 -920
<< locali >>
rect 240 -1020 450 -920
use n1x30  n1x30_0
timestamp 1732727030
transform 1 0 -180 0 1 -120
box -500 -1000 600 300
use n1x30  n1x30_2
timestamp 1732727030
transform -1 0 850 0 1 -120
box -500 -1000 600 300
<< labels >>
flabel space -100 30 -100 30 0 FreeSans 800 0 0 0 DL
port 0 nsew
flabel space 760 30 760 30 0 FreeSans 800 0 0 0 DR
port 1 nsew
flabel space -580 -470 -580 -470 0 FreeSans 800 0 0 0 GL
port 2 nsew
flabel space 1250 -480 1250 -480 0 FreeSans 800 0 0 0 GR
port 3 nsew
flabel space -90 -970 -90 -970 0 FreeSans 800 0 0 0 S
port 4 nsew
flabel space -580 80 -580 80 0 FreeSans 800 0 0 0 B
port 5 nsew
<< end >>
