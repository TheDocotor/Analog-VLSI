magic
tech sky130A
magscale 1 2
timestamp 1730763487
<< nwell >>
rect 150 1547 2950 1550
rect 134 -468 2965 1547
<< nsubdiff >>
rect 173 1495 2926 1508
rect 173 -403 199 1495
rect 238 1430 2861 1456
rect 238 -351 251 1430
rect 2848 -264 2861 1430
rect 2848 -351 2861 -303
rect 238 -364 2861 -351
rect 2900 -403 2926 1495
rect 173 -429 2926 -403
<< nsubdiffcont >>
rect 199 1456 2900 1495
rect 199 -364 238 1456
rect 2861 -264 2900 1456
rect 2848 -303 2900 -264
rect 2861 -364 2900 -303
rect 199 -403 2900 -364
<< locali >>
rect 173 1495 2926 1508
rect 173 -403 199 1495
rect 238 1430 2861 1456
rect 238 -351 251 1430
rect 2848 -264 2861 1430
rect 2848 -351 2861 -303
rect 238 -364 2861 -351
rect 2900 -403 2926 1495
rect 173 -429 2926 -403
<< viali >>
rect 750 -225 1300 -175
rect 1600 -225 2150 -175
rect 750 -675 1300 -625
rect 1600 -675 2150 -625
<< metal1 >>
rect 725 -175 1325 -150
rect 725 -225 750 -175
rect 1300 -225 1325 -175
rect 725 -625 1325 -225
rect 725 -675 750 -625
rect 1300 -675 1325 -625
rect 725 -700 1325 -675
rect 1575 -175 2175 -150
rect 1575 -225 1600 -175
rect 2150 -225 2175 -175
rect 1575 -625 2175 -225
rect 1575 -675 1600 -625
rect 2150 -675 2175 -625
rect 1575 -700 2175 -675
use n20x1  n20x1_1
timestamp 1730763316
transform -1 0 2600 0 1 -1100
box -300 -1200 1200 600
use n20x1  n20x1_2
timestamp 1730763316
transform 1 0 550 0 1 -1100
box -300 -1200 1200 600
use p20x1  p20x1_0
timestamp 1730763316
transform 1 0 525 0 -1 250
box -225 -1150 1075 550
use p20x1  p20x1_1
timestamp 1730763316
transform -1 0 2575 0 -1 250
box -225 -1150 1075 550
<< end >>
