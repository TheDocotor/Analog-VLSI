magic
tech sky130A
timestamp 1731631080
<< xpolycontact >>
rect -142 -609 -107 -393
rect 107 -609 142 -393
<< xpolyres >>
rect -142 574 -24 609
rect -142 -393 -107 574
rect -59 -306 -24 574
rect 24 574 142 609
rect 24 -306 59 574
rect -59 -341 59 -306
rect 107 -393 142 574
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 9.5 m 1 nx 4 wmin 0.350 lmin 0.50 rho 2000 val 224.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_0p35_FNGBKB parameters
<< end >>
