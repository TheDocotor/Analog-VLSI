magic
tech sky130A
magscale 1 2
timestamp 1730605901
<< xpolycontact >>
rect -573 16452 573 16884
rect -573 52 573 484
rect -573 -484 573 -52
rect -573 -16884 573 -16452
<< xpolyres >>
rect -573 484 573 16452
rect -573 -16452 573 -484
<< viali >>
rect -557 16469 557 16866
rect -557 70 557 467
rect -557 -467 557 -70
rect -557 -16866 557 -16469
<< metal1 >>
rect -569 16866 569 16872
rect -569 16469 -557 16866
rect 557 16469 569 16866
rect -569 16463 569 16469
rect -569 467 569 473
rect -569 70 -557 467
rect 557 70 569 467
rect -569 64 569 70
rect -569 -70 569 -64
rect -569 -467 -557 -70
rect 557 -467 569 -70
rect -569 -473 569 -467
rect -569 -16469 569 -16463
rect -569 -16866 -557 -16469
rect 557 -16866 569 -16469
rect -569 -16872 569 -16866
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 80 m 2 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 27.988k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_5p73_YK3U8H parameters
<< end >>
