magic
tech sky130A
magscale 1 2
timestamp 1732920865
<< nwell >>
rect -2200 5359 6000 5360
rect -2202 4400 6000 5359
rect 1110 3750 1280 3790
rect 4080 3740 6000 4400
<< pwell >>
rect -6800 5400 13400 8100
rect -6800 4370 -2250 5400
rect -6800 3850 4020 4370
rect -6800 3847 -84 3850
rect 2716 3847 4020 3850
rect -6800 1832 -100 3847
rect 2731 3720 4020 3847
rect 6160 4370 13400 5400
rect 6070 3720 13400 4370
rect 2731 1832 13400 3720
rect -6800 -10500 13400 1832
rect -6800 -16860 3800 -10500
rect -6800 -16900 10180 -16860
rect 10200 -16900 13400 -10500
rect -6800 -18000 13400 -16900
<< pmos >>
rect -1500 4694 -1300 4894
rect -1180 4694 -980 4894
<< pdiff >>
rect -1500 4940 -1300 4952
rect -1500 4906 -1488 4940
rect -1312 4906 -1300 4940
rect -1500 4894 -1300 4906
rect -1180 4940 -980 4952
rect -1180 4906 -1168 4940
rect -992 4906 -980 4940
rect -1180 4894 -980 4906
rect -1500 4682 -1300 4694
rect -1500 4648 -1488 4682
rect -1312 4648 -1300 4682
rect -1500 4636 -1300 4648
rect -1180 4682 -980 4694
rect -1180 4648 -1168 4682
rect -992 4648 -980 4682
rect -1180 4636 -980 4648
<< pdiffc >>
rect -1488 4906 -1312 4940
rect -1168 4906 -992 4940
rect -1488 4648 -1312 4682
rect -1168 4648 -992 4682
<< psubdiff >>
rect -6800 7900 13400 8100
rect -6800 7500 -6400 7900
rect 13000 7500 13400 7900
rect -6800 7300 13400 7500
rect -6800 5200 -6000 7300
rect 12600 5400 13400 7300
rect -6800 -17000 -6600 5200
rect -6200 -17000 -6000 5200
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect -6800 -17200 -6000 -17000
rect 12600 -17200 13400 -16800
rect -6800 -17400 13400 -17200
rect -6800 -17800 -6200 -17400
rect 13000 -17800 13400 -17400
rect -6800 -18000 13400 -17800
<< nsubdiff >>
rect -2110 5275 5920 5300
rect -2110 5180 -2075 5275
rect -2100 4525 -2075 5180
rect -2025 5260 5920 5275
rect -2025 5220 -1880 5260
rect 5740 5220 5920 5260
rect -2025 5180 5920 5220
rect -2025 4575 -2000 5180
rect 5840 5120 5920 5180
rect -2025 4540 4250 4575
rect -2025 4525 -1970 4540
rect -2100 4500 -1970 4525
rect 4180 4500 4250 4540
rect -2100 4480 4250 4500
rect 4160 4475 4250 4480
rect 4160 4460 4240 4475
rect 4160 3880 4180 4460
rect 4220 3900 4240 4460
rect 5840 3960 5860 5120
rect 5900 3960 5920 5120
rect 5840 3900 5920 3960
rect 4220 3880 5920 3900
rect 4160 3840 4270 3880
rect 5840 3840 5920 3880
rect 4160 3820 5920 3840
<< psubdiffcont >>
rect -6400 7500 13000 7900
rect -6600 -17000 -6200 5200
rect 12800 -16800 13200 5400
rect -6200 -17800 13000 -17400
<< nsubdiffcont >>
rect -2075 4525 -2025 5275
rect -1880 5220 5740 5260
rect -1970 4500 4180 4540
rect 4180 3880 4220 4460
rect 5860 3960 5900 5120
rect 4270 3840 5840 3880
<< poly >>
rect -1597 4878 -1500 4894
rect -1597 4710 -1581 4878
rect -1547 4710 -1500 4878
rect -1597 4694 -1500 4710
rect -1300 4694 -1180 4894
rect -980 4878 -883 4894
rect -980 4710 -933 4878
rect -899 4710 -883 4878
rect -980 4694 -883 4710
rect -2310 4250 -2254 4258
rect -2380 4220 -2254 4250
rect -2380 4100 -2360 4220
rect -2300 4100 -2254 4220
rect -2380 4060 -2254 4100
rect -2310 4058 -2254 4060
rect -1740 3180 -1710 3250
rect -1750 3160 -1640 3180
rect -1750 3060 -1700 3160
rect -1660 3060 -1640 3160
rect -1750 3050 -1640 3060
rect -1740 3040 -1640 3050
rect -1740 -16810 -1710 3040
rect -280 1180 -220 1280
<< polycont >>
rect -1581 4710 -1547 4878
rect -933 4710 -899 4878
rect -2360 4100 -2300 4220
rect -1700 3060 -1660 3160
<< locali >>
rect -6800 7900 13400 8100
rect -6800 7500 -6400 7900
rect 13000 7500 13400 7900
rect -6800 7300 13400 7500
rect -6800 5200 -3800 7300
rect 12600 5400 13400 7300
rect -6800 -17000 -6600 5200
rect -6200 3200 -3800 5200
rect -2110 5275 5920 5300
rect -2110 5180 -2075 5275
rect -2100 4525 -2075 5180
rect -2025 5260 5920 5275
rect -2025 5220 -1880 5260
rect 5740 5220 5920 5260
rect -2025 5180 5920 5220
rect -2025 4575 -2000 5180
rect 5840 5120 5920 5180
rect -1504 4906 -1488 4940
rect -1312 4906 -1296 4940
rect -1184 4906 -1168 4940
rect -992 4906 -976 4940
rect -1581 4878 -1547 4894
rect -933 4878 -899 4894
rect -1547 4710 -1540 4720
rect -1581 4700 -1540 4710
rect -1581 4694 -1500 4700
rect -933 4694 -899 4710
rect -1580 4682 -1500 4694
rect -1580 4648 -1488 4682
rect -1312 4648 -1296 4682
rect -1184 4648 -1168 4682
rect -992 4648 -976 4682
rect -1580 4640 -1500 4648
rect -2025 4540 4250 4575
rect -2025 4525 -1970 4540
rect -2100 4500 -1970 4525
rect 4180 4500 4250 4540
rect -2100 4480 4250 4500
rect 4160 4475 4250 4480
rect 4160 4460 4240 4475
rect -2370 4220 -2290 4240
rect -2370 4100 -2360 4220
rect -2300 4100 -2290 4220
rect -2370 4080 -2290 4100
rect 4160 3880 4180 4460
rect 4220 3900 4240 4460
rect 5840 3960 5860 5120
rect 5900 3960 5920 5120
rect 5840 3900 5920 3960
rect 4220 3880 5920 3900
rect 4160 3840 4270 3880
rect 5840 3840 5920 3880
rect 4160 3820 5920 3840
rect -6200 -2042 -6000 3200
rect -1720 3160 -1640 3180
rect -1720 3060 -1700 3160
rect -1660 3060 -1640 3160
rect -1720 3040 -1640 3060
rect 2320 1420 2570 1700
rect 480 -60 1960 140
rect -1440 -460 1960 -60
rect -6200 -17000 -6009 -2042
rect -5000 -13200 -2200 -12800
rect -6800 -17209 -6009 -17000
rect -1840 -16822 -1760 -16820
rect -1840 -16856 -1832 -16822
rect -1772 -16856 -1760 -16822
rect -1840 -17200 -1760 -16856
rect -1000 -17200 1200 -460
rect 3740 -10660 10180 -10440
rect 3740 -11500 3960 -10660
rect 4800 -11500 5240 -10660
rect 6100 -11500 6540 -10660
rect 7380 -11500 7820 -10660
rect 8680 -11500 9120 -10660
rect 9940 -11500 10160 -10660
rect 3740 -11940 10180 -11500
rect 3740 -12780 3960 -11940
rect 4800 -12780 5240 -11940
rect 6100 -12780 6540 -11940
rect 7380 -12780 7820 -11940
rect 8680 -12780 9120 -11940
rect 9940 -12780 10160 -11940
rect 3740 -13220 10180 -12780
rect 3740 -14080 3960 -13220
rect 4800 -14080 5240 -13220
rect 6100 -14080 6540 -13220
rect 7380 -14080 7820 -13220
rect 8680 -14080 9120 -13220
rect 9940 -14080 10160 -13220
rect 3740 -14520 10180 -14080
rect 3740 -15360 3960 -14520
rect 4800 -15360 5240 -14520
rect 6100 -15360 6540 -14520
rect 7380 -15360 7820 -14520
rect 8680 -15360 9120 -14520
rect 9940 -15360 10160 -14520
rect 3740 -15800 10180 -15360
rect 3740 -16640 3960 -15800
rect 4800 -16640 5240 -15800
rect 6100 -16640 6540 -15800
rect 7380 -16640 7820 -15800
rect 8680 -16640 9120 -15800
rect 9940 -16640 10160 -15800
rect 3740 -16940 10180 -16640
rect 3340 -17200 10180 -16940
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect 12600 -17200 13400 -16800
rect -2203 -17209 13400 -17200
rect -6800 -17400 13400 -17209
rect -6800 -17800 -6200 -17400
rect 13000 -17800 13400 -17400
rect -6800 -18000 13400 -17800
<< viali >>
rect -6400 7500 13000 7900
rect 6720 6220 7500 6440
rect 8340 6200 9020 6440
rect -6600 -17000 -6200 5200
rect -2075 4525 -2025 5275
rect -1880 5220 5740 5260
rect 4750 4995 5500 5045
rect -1488 4906 -1312 4940
rect -1168 4906 -992 4940
rect 1112 4906 1288 4940
rect -1581 4710 -1547 4878
rect -933 4710 -899 4878
rect 1019 4710 1053 4878
rect -1488 4648 -1312 4682
rect -1168 4648 -992 4682
rect 1112 4648 1288 4682
rect -1970 4500 4180 4540
rect 1120 4400 1280 4440
rect -1500 4270 -1300 4304
rect -1140 4280 -1000 4340
rect -2360 4100 -2300 4220
rect -2242 4012 -1266 4046
rect 4180 3880 4220 4460
rect 4360 4280 4400 4340
rect 4750 3995 5500 4045
rect 5860 3960 5900 5120
rect 4270 3840 5840 3880
rect 1832 3756 2002 3796
rect -3412 3307 -2298 3704
rect 1120 3600 1280 3640
rect -1832 3260 -1772 3294
rect -1700 3060 -1660 3160
rect -1175 3025 -625 3075
rect -280 2850 -220 2950
rect 2480 2540 2540 2740
rect 120 2220 160 2320
rect -280 1180 -220 1280
rect 140 800 180 1000
rect 2500 800 2540 1000
rect -1832 -16856 -1772 -16822
rect 1776 -9743 2890 -9346
rect 6940 -10180 7300 -9980
rect 8600 -10200 8760 -9960
rect 1776 -14142 2890 -13745
rect 12800 -16800 13200 5400
rect -6200 -17800 13000 -17400
<< metal1 >>
rect -6800 7900 13400 8100
rect -6800 7500 -6400 7900
rect 13000 7500 13400 7900
rect -6800 7300 13400 7500
rect -6800 5200 -3800 7300
rect 6680 6440 7540 6460
rect 6680 6220 6720 6440
rect 7500 6220 7540 6440
rect 6680 6180 7540 6220
rect 8320 6440 9040 6460
rect 8320 6200 8340 6440
rect 9020 6200 9040 6440
rect 8320 6180 9040 6200
rect -6800 -17000 -6600 5200
rect -6200 3200 -3800 5200
rect -2200 5275 6000 5640
rect -2200 5120 -2075 5275
rect -2120 4525 -2075 5120
rect -2025 5260 6000 5275
rect -2025 5220 -1880 5260
rect 5740 5220 6000 5260
rect -2025 5120 6000 5220
rect 12600 5400 13400 7300
rect -2025 4575 -2000 5120
rect -1500 4940 -1300 5120
rect -1500 4906 -1488 4940
rect -1312 4906 -1300 4940
rect -1500 4900 -1300 4906
rect -1180 4940 -980 5120
rect -1180 4906 -1168 4940
rect -992 4906 -980 4940
rect -1180 4900 -980 4906
rect 1100 4940 1300 5120
rect 4740 5045 5530 5120
rect 4740 4995 4750 5045
rect 5500 4995 5530 5045
rect 4740 4980 5530 4995
rect 1100 4906 1112 4940
rect 1288 4906 1300 4940
rect 1100 4900 1300 4906
rect -1587 4878 -1541 4890
rect -939 4880 -893 4890
rect -1587 4710 -1581 4878
rect -1547 4710 -1541 4878
rect -1587 4698 -1541 4710
rect -940 4878 1060 4880
rect -940 4710 -933 4878
rect -899 4710 1019 4878
rect 1053 4710 1060 4878
rect -940 4700 1060 4710
rect -939 4698 -893 4700
rect -1500 4682 -1300 4688
rect -1500 4630 -1490 4682
rect -1310 4630 -1300 4682
rect -1500 4620 -1300 4630
rect -1180 4682 -980 4688
rect -1180 4630 -1170 4682
rect -990 4630 -980 4682
rect -1180 4620 -980 4630
rect 1100 4630 1110 4680
rect 1290 4630 1300 4680
rect 1100 4620 1300 4630
rect -2025 4540 4250 4575
rect -2025 4525 -1970 4540
rect -2120 4500 -1970 4525
rect 4180 4500 4250 4540
rect -2120 4480 4250 4500
rect 4160 4475 4250 4480
rect 4160 4460 4240 4475
rect 1100 4442 1300 4450
rect 1100 4390 1120 4442
rect 1280 4390 1300 4442
rect -1180 4340 -980 4350
rect -1510 4330 -1290 4340
rect -1510 4320 -1500 4330
rect -1520 4270 -1500 4320
rect -1300 4320 -1290 4330
rect -1300 4270 -1280 4320
rect -1520 4260 -1280 4270
rect -1180 4280 -1140 4340
rect -1000 4280 -980 4340
rect -2380 4220 -2280 4240
rect -2380 4100 -2360 4220
rect -2300 4100 -2280 4220
rect -2380 4080 -2280 4100
rect -2255 4050 -1255 4055
rect -2260 4046 -1240 4050
rect -2260 4040 -2242 4046
rect -2620 4012 -2242 4040
rect -1266 4012 -1240 4046
rect -2620 3852 -1240 4012
rect -3332 3722 -1240 3852
rect -3428 3704 -1240 3722
rect -3428 3307 -3412 3704
rect -2298 3500 -1240 3704
rect -2298 3420 -2186 3500
rect -2298 3307 -2282 3420
rect -3428 3290 -2282 3307
rect -1180 3300 -980 4280
rect 1100 3810 1300 4390
rect 4160 3880 4180 4460
rect 4220 3900 4240 4460
rect 4340 4340 4420 4360
rect 4400 4280 4420 4340
rect 4340 4260 4420 4280
rect 4720 4050 5520 4060
rect 4720 3995 4750 4050
rect 5500 3995 5520 4050
rect 4720 3980 5520 3995
rect 5840 3960 5860 5120
rect 5900 3960 5920 5120
rect 5840 3900 5920 3960
rect 4220 3880 5920 3900
rect 4160 3840 4270 3880
rect 5840 3840 5920 3880
rect 4160 3820 5920 3840
rect 1100 3796 2030 3810
rect 1100 3756 1832 3796
rect 2002 3756 2030 3796
rect 1100 3730 2030 3756
rect 1100 3640 1300 3730
rect 1100 3600 1120 3640
rect 1280 3600 1300 3640
rect 1100 3580 1300 3600
rect -1840 3294 -980 3300
rect -1840 3260 -1832 3294
rect -1772 3260 -980 3294
rect -6200 -2042 -6000 3200
rect -1655 3185 -1610 3260
rect -1700 3170 -1610 3185
rect -1720 3160 -1610 3170
rect -1720 3060 -1700 3160
rect -1660 3155 -1610 3160
rect -1660 3060 -1650 3155
rect -1180 3140 -980 3260
rect -1180 3100 -600 3140
rect -1720 3050 -1650 3060
rect -1710 3040 -1650 3050
rect -1200 3075 -600 3100
rect -1200 3025 -1175 3075
rect -625 3025 -600 3075
rect -1200 3000 -600 3025
rect -300 2950 -200 2970
rect -300 2850 -280 2950
rect -220 2850 -200 2950
rect -300 2830 -200 2850
rect 2460 2740 2560 2760
rect 2460 2540 2480 2740
rect 2540 2540 2560 2740
rect 2460 2520 2560 2540
rect 100 2320 180 2340
rect 100 2220 120 2320
rect 100 2200 180 2220
rect -200 1700 500 1800
rect -200 1300 -60 1700
rect -300 1280 -60 1300
rect -300 1180 -280 1280
rect -220 1180 -60 1280
rect -300 1160 -60 1180
rect 120 1000 200 1020
rect 120 800 140 1000
rect 120 780 200 800
rect 2480 1000 2560 1020
rect 2540 800 2560 1000
rect 2480 780 2560 800
rect 480 -60 1960 140
rect -1440 -460 1960 -60
rect -6200 -17000 -6009 -2042
rect -5000 -13200 -2200 -12800
rect -6800 -17209 -6009 -17000
rect -1840 -16822 -1760 -16820
rect -1840 -16856 -1832 -16822
rect -1772 -16856 -1760 -16822
rect -1840 -17200 -1760 -16856
rect -1000 -17200 1200 -460
rect 1740 -9346 2620 -9320
rect 2800 -9346 6020 -9320
rect 1740 -9743 1776 -9346
rect 2890 -9743 6020 -9346
rect 1740 -9760 2620 -9743
rect 2800 -9760 6020 -9743
rect 5440 -9880 6020 -9760
rect 5440 -9980 7740 -9880
rect 5440 -10180 6940 -9980
rect 7300 -10180 7740 -9980
rect 5440 -10300 7740 -10180
rect 8540 -9960 8840 -9940
rect 8540 -10200 8600 -9960
rect 8760 -10200 8840 -9960
rect 8540 -10260 8840 -10200
rect 4080 -11380 9860 -10760
rect 4080 -12060 4700 -11380
rect 5360 -12060 5980 -11380
rect 6660 -12060 7260 -11380
rect 7940 -12060 8560 -11380
rect 9240 -12060 9860 -11380
rect 4080 -12680 9860 -12060
rect 4080 -13730 4700 -12680
rect 1760 -13745 4700 -13730
rect 1760 -14142 1776 -13745
rect 2890 -14142 4700 -13745
rect 1760 -14160 4700 -14142
rect 4080 -14640 4700 -14160
rect 5360 -14640 5980 -12680
rect 7940 -14640 8560 -12680
rect 9240 -14640 9860 -12680
rect 4080 -15260 9860 -14640
rect 4080 -15920 4700 -15260
rect 5360 -15920 5980 -15260
rect 6660 -15920 7260 -15260
rect 7940 -15920 8560 -15260
rect 9240 -15920 9860 -15260
rect 4080 -16540 9860 -15920
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect 3740 -16940 10180 -16860
rect 3340 -17200 10180 -16940
rect 12600 -17200 13400 -16800
rect -2203 -17209 13400 -17200
rect -6800 -17400 13400 -17209
rect -6800 -17800 -6200 -17400
rect 13000 -17800 13400 -17400
rect -6800 -18000 13400 -17800
<< via1 >>
rect 6720 6220 7500 6440
rect 8340 6200 9020 6440
rect -1490 4648 -1488 4682
rect -1488 4648 -1312 4682
rect -1312 4648 -1310 4682
rect -1490 4630 -1310 4648
rect -1170 4648 -1168 4682
rect -1168 4648 -992 4682
rect -992 4648 -990 4682
rect -1170 4630 -990 4648
rect 1110 4648 1112 4682
rect 1112 4648 1288 4682
rect 1288 4648 1290 4682
rect 1110 4630 1290 4648
rect 1120 4440 1280 4442
rect 1120 4400 1280 4440
rect 1120 4390 1280 4400
rect -1500 4304 -1300 4330
rect -1500 4270 -1300 4304
rect -1140 4280 -1000 4340
rect -2360 4100 -2300 4220
rect 4340 4280 4360 4340
rect 4360 4280 4400 4340
rect 4750 4045 5500 4050
rect 4750 3995 5500 4045
rect -280 2850 -220 2950
rect 2480 2540 2540 2740
rect 120 2220 160 2320
rect 160 2220 180 2320
rect 140 800 180 1000
rect 180 800 200 1000
rect 2480 800 2500 1000
rect 2500 800 2540 1000
rect 1776 -9743 2890 -9346
rect 8600 -10200 8760 -9960
rect 6740 -13800 7150 -13530
<< metal2 >>
rect 6360 6520 6500 6540
rect 6360 6440 9240 6520
rect 6360 6220 6720 6440
rect 7500 6220 8340 6440
rect 6360 6200 8340 6220
rect 9020 6200 9240 6440
rect 6360 6120 9240 6200
rect -1500 4682 -1300 4690
rect -1500 4630 -1490 4682
rect -1310 4630 -1300 4682
rect -1500 4340 -1300 4630
rect -1180 4682 -980 4690
rect -1180 4630 -1170 4682
rect -990 4630 -980 4682
rect -1180 4360 -980 4630
rect 1100 4682 1300 4690
rect 1100 4630 1110 4682
rect 1290 4630 1300 4682
rect 1100 4442 1300 4630
rect 1100 4390 1120 4442
rect 1280 4390 1300 4442
rect -1180 4340 4400 4360
rect -1520 4330 -1280 4340
rect -1520 4270 -1500 4330
rect -1300 4270 -1280 4330
rect -1520 4260 -1280 4270
rect -1180 4280 -1140 4340
rect -1000 4280 4340 4340
rect -1180 4260 4400 4280
rect -2380 4220 -2280 4240
rect -2380 4100 -2360 4220
rect -2300 4205 -2255 4220
rect -2300 4200 -480 4205
rect -2300 4140 3680 4200
rect -2300 4125 -2255 4140
rect -2300 4100 -2280 4125
rect -2380 4080 -2280 4100
rect -420 4080 3680 4140
rect -280 2970 -230 4080
rect 3540 3770 3680 4080
rect 4720 4050 5520 4060
rect 4720 3995 4750 4050
rect 5500 3995 5520 4050
rect 4720 3780 5520 3995
rect 6360 3780 6500 6120
rect 4720 3770 6500 3780
rect 3540 3670 6500 3770
rect 5400 3660 6500 3670
rect -300 2950 -200 2970
rect -300 2850 -280 2950
rect -220 2850 -200 2950
rect -300 2830 -200 2850
rect 2460 2740 4380 2760
rect 2460 2540 2480 2740
rect 2540 2540 4380 2740
rect 2460 2520 4380 2540
rect 100 2320 2860 2340
rect 100 2220 120 2320
rect 180 2220 2860 2320
rect 100 2200 2860 2220
rect 100 1000 2560 1020
rect 100 800 140 1000
rect 200 800 2480 1000
rect 2540 800 2560 1000
rect 100 780 2560 800
rect 2700 -8780 2860 2200
rect 3940 -1800 4380 2520
rect 3940 -2140 9000 -1800
rect 2540 -9320 2860 -8780
rect 1740 -9346 2900 -9320
rect 1740 -9743 1776 -9346
rect 2890 -9743 2900 -9346
rect 1740 -9760 2900 -9743
rect 8500 -9960 9000 -2140
rect 8500 -10200 8600 -9960
rect 8760 -10200 9000 -9960
rect 8500 -13400 9000 -10200
rect 6700 -13530 9000 -13400
rect 6700 -13800 6740 -13530
rect 7150 -13800 9000 -13530
rect 6700 -13900 9000 -13800
use diff_pair  diff_pair_0
timestamp 1730763487
transform 1 0 -234 0 1 2300
box 134 -2300 2965 1550
use n20x1  n20x1_0
timestamp 1730763316
transform -1 0 -400 0 1 2600
box -300 -1200 1200 600
use n20x1  n20x1_1
timestamp 1730763316
transform -1 0 -400 0 1 1000
box -300 -1200 1200 600
use p20x05  p20x05_0
timestamp 1730605901
transform 1 0 1825 0 1 3470
box 2475 450 3975 1650
use sky130_fd_pr__nfet_01v8_6EEDFX  sky130_fd_pr__nfet_01v8_6EEDFX_0
timestamp 1730747568
transform 0 1 -1754 -1 0 4158
box -158 -526 158 526
use sky130_fd_pr__nfet_01v8_N7YW8T  sky130_fd_pr__nfet_01v8_N7YW8T_0
timestamp 1730605901
transform 0 1 -1802 -1 0 -1752
box -5058 -68 5058 68
use sky130_fd_pr__nfet_01v8_N7YW8T  sky130_fd_pr__nfet_01v8_N7YW8T_1
timestamp 1730605901
transform 0 1 -1802 -1 0 -11810
box -5058 -68 5058 68
use sky130_fd_pr__pfet_01v8_J24L55  sky130_fd_pr__pfet_01v8_J24L55_0
timestamp 1730316371
transform 0 1 1200 -1 0 4794
box -194 -200 194 200
use sky130_fd_pr__res_xhigh_po_5p73_G7V36E  sky130_fd_pr__res_xhigh_po_5p73_G7V36E_0
timestamp 1730769459
transform 1 0 2333 0 1 -11744
box -573 -2416 573 2416
use sky130_fd_pr__res_xhigh_po_5p73_J2M2GK  sky130_fd_pr__res_xhigh_po_5p73_J2M2GK_0
timestamp 1730769459
transform 1 0 -2855 0 1 -4694
box -573 -8416 573 8416
use sky130_fd_pr__res_xhigh_po_5p73_J2M2GK  sky130_fd_pr__res_xhigh_po_5p73_J2M2GK_1
timestamp 1730769459
transform 1 0 -4427 0 1 -4784
box -573 -8416 573 8416
use sky130_fd_pr__res_xhigh_po_5p73_J2MYFK  sky130_fd_pr__res_xhigh_po_5p73_J2MYFK_0
timestamp 1730769459
transform 1 0 7173 0 1 -1884
box -573 -8416 573 8416
use sky130_fd_pr__res_xhigh_po_5p73_J2MYFK  sky130_fd_pr__res_xhigh_po_5p73_J2MYFK_1
timestamp 1730769459
transform 1 0 8673 0 1 -1884
box -573 -8416 573 8416
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 4 1288
timestamp 1704896540
transform 1 0 3716 0 1 -16896
box 0 0 1340 1340
<< labels >>
flabel metal1 200 5400 200 5400 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 1220 3980 1220 3980 0 FreeSans 800 0 0 0 Vdiff
flabel metal1 -1840 3730 -1840 3730 0 FreeSans 800 0 0 0 Vres
flabel metal1 -1090 3730 -1090 3730 0 FreeSans 800 0 0 0 Vdm2
flabel viali 1030 4800 1030 4800 0 FreeSans 800 0 0 0 Vpgates
flabel metal2 2720 -9340 2720 -9340 0 FreeSans 800 0 0 0 diffg1
flabel metal2 5700 3700 5700 3700 0 FreeSans 1600 0 0 0 Vref
port 1 nsew
flabel metal1 -6460 -17640 -6460 -17640 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
<< end >>
