magic
tech sky130A
magscale 1 2
timestamp 1730605901
<< nwell >>
rect -2200 5359 6000 5360
rect -2202 4400 6000 5359
rect 4080 3740 6000 4400
<< pwell >>
rect -9800 5360 13400 6800
rect -9800 5359 -2200 5360
rect -9800 4400 -2202 5359
rect -9800 3850 4080 4400
rect -9800 3847 16 3850
rect 2416 3847 4080 3850
rect -9800 1832 0 3847
rect 2431 3740 4080 3847
rect 6000 3740 13400 5360
rect 2431 1832 13400 3740
rect -9800 -3400 13400 1832
rect -9800 -9760 3800 -3400
rect -9800 -9800 10180 -9760
rect 10200 -9800 13400 -3400
rect -9800 -18000 13400 -9800
<< pmos >>
rect -1500 4694 -1300 4894
rect -1180 4694 -980 4894
<< pdiff >>
rect -1500 4940 -1300 4952
rect -1500 4906 -1488 4940
rect -1312 4906 -1300 4940
rect -1500 4894 -1300 4906
rect -1180 4940 -980 4952
rect -1180 4906 -1168 4940
rect -992 4906 -980 4940
rect -1180 4894 -980 4906
rect -1500 4682 -1300 4694
rect -1500 4648 -1488 4682
rect -1312 4648 -1300 4682
rect -1500 4636 -1300 4648
rect -1180 4682 -980 4694
rect -1180 4648 -1168 4682
rect -992 4648 -980 4682
rect -1180 4636 -980 4648
<< pdiffc >>
rect -1488 4906 -1312 4940
rect -1168 4906 -992 4940
rect -1488 4648 -1312 4682
rect -1168 4648 -992 4682
<< psubdiff >>
rect -9800 6600 13400 6800
rect -9800 6200 -9400 6600
rect 13000 6200 13400 6600
rect -9800 6000 13400 6200
rect -9800 5200 -9000 6000
rect 12600 5400 13400 6000
rect -9800 -17000 -9600 5200
rect -9200 -17000 -9000 5200
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect -9800 -17200 -9000 -17000
rect 12600 -17200 13400 -16800
rect -9800 -17400 13400 -17200
rect -9800 -17800 -9200 -17400
rect 13000 -17800 13400 -17400
rect -9800 -18000 13400 -17800
<< mvnsubdiff >>
rect -2120 5260 5920 5280
rect -2120 5240 -2020 5260
rect -2120 4520 -2100 5240
rect -2060 5220 -2020 5240
rect 5860 5220 5920 5260
rect -2060 5180 5920 5220
rect -2060 4560 -2040 5180
rect -2060 4540 4240 4560
rect -2060 4520 -2020 4540
rect -2120 4500 -2020 4520
rect 4160 4500 4240 4540
rect -2120 4480 4240 4500
rect 4160 4420 4240 4480
rect 4160 3940 4180 4420
rect 4220 3940 4240 4420
rect 4160 3900 4240 3940
rect 5840 3920 5860 5180
rect 5900 3920 5920 5180
rect 5840 3900 5920 3920
rect 4160 3880 5920 3900
rect 4160 3840 4200 3880
rect 5820 3840 5920 3880
rect 4160 3820 5920 3840
<< psubdiffcont >>
rect -9400 6200 13000 6600
rect -9600 -17000 -9200 5200
rect 12800 -16800 13200 5400
rect -9200 -17800 13000 -17400
<< mvnsubdiffcont >>
rect -2100 4520 -2060 5240
rect -2020 5220 5860 5260
rect -2020 4500 4160 4540
rect 4180 3940 4220 4420
rect 5860 3920 5900 5180
rect 4200 3840 5820 3880
<< poly >>
rect -1597 4878 -1500 4894
rect -1597 4710 -1581 4878
rect -1547 4710 -1500 4878
rect -1597 4694 -1500 4710
rect -1300 4694 -1180 4894
rect -980 4878 -883 4894
rect -980 4710 -933 4878
rect -899 4710 -883 4878
rect -980 4694 -883 4710
rect -2310 4058 -2254 4258
rect -1750 3055 -1745 3170
rect -1740 -16810 -1710 3250
<< polycont >>
rect -1581 4710 -1547 4878
rect -933 4710 -899 4878
<< locali >>
rect -9800 6600 13400 6800
rect -9800 6200 -9400 6600
rect 13000 6200 13400 6600
rect -9800 6000 13400 6200
rect -9800 5200 -9000 6000
rect 12600 5400 13400 6000
rect -9800 -17000 -9600 5200
rect -9200 -2080 -9000 5200
rect -2120 5260 5920 5280
rect -2120 5240 -2020 5260
rect -2120 4520 -2100 5240
rect -2060 5220 -2020 5240
rect 5860 5220 5920 5260
rect -2060 5180 5920 5220
rect -2060 4560 -2040 5180
rect -1504 4906 -1488 4940
rect -1312 4906 -1296 4940
rect -1184 4906 -1168 4940
rect -992 4906 -976 4940
rect -1581 4878 -1547 4894
rect -933 4878 -899 4894
rect -1547 4710 -1540 4720
rect -1581 4700 -1540 4710
rect -1581 4694 -1500 4700
rect -933 4694 -899 4710
rect -1580 4682 -1500 4694
rect -1580 4648 -1488 4682
rect -1312 4648 -1296 4682
rect -1184 4648 -1168 4682
rect -992 4648 -976 4682
rect -1580 4640 -1500 4648
rect -2060 4540 4240 4560
rect -2060 4520 -2020 4540
rect -2120 4500 -2020 4520
rect 4160 4500 4240 4540
rect -2120 4480 4240 4500
rect 4160 4420 4240 4480
rect 4160 3940 4180 4420
rect 4220 3940 4240 4420
rect 4160 3900 4240 3940
rect 5840 3920 5860 5180
rect 5900 3920 5920 5180
rect 5840 3900 5920 3920
rect 4160 3880 5920 3900
rect 4160 3840 4200 3880
rect 5820 3840 5920 3880
rect 4160 3820 5920 3840
rect 5520 3460 5840 3480
rect -1750 3170 -1715 3180
rect -1750 3050 -1715 3055
rect 5790 2690 5840 3460
rect 5520 2560 5840 2690
rect 2020 1000 2180 1580
rect 2020 800 2160 1000
rect 2020 420 2180 800
rect 480 -60 1960 140
rect -1440 -460 1960 -60
rect -9200 -17000 -2180 -2080
rect -9800 -17200 -2180 -17000
rect -1840 -16822 -1760 -16820
rect -1840 -16856 -1832 -16822
rect -1772 -16856 -1760 -16822
rect -1840 -17200 -1760 -16856
rect -1000 -17200 1200 -460
rect 1760 -1620 2880 -1360
rect 1760 -2100 2640 -1620
rect 2780 -2100 2880 -1620
rect 1760 -2660 2880 -2100
rect 3740 -3560 10180 -3340
rect 3740 -4400 3960 -3560
rect 4800 -4400 5240 -3560
rect 6100 -4400 6540 -3560
rect 7380 -4400 7820 -3560
rect 8680 -4400 9120 -3560
rect 9940 -4400 10160 -3560
rect 3740 -4840 10180 -4400
rect 3740 -5680 3960 -4840
rect 4800 -5680 5240 -4840
rect 6100 -5680 6540 -4840
rect 7380 -5680 7820 -4840
rect 8680 -5680 9120 -4840
rect 9940 -5680 10160 -4840
rect 3740 -6120 10180 -5680
rect 3740 -6980 3960 -6120
rect 4800 -6980 5240 -6120
rect 6100 -6980 6540 -6120
rect 7380 -6980 7820 -6120
rect 8680 -6980 9120 -6120
rect 9940 -6980 10160 -6120
rect 3740 -7420 10180 -6980
rect 3740 -8260 3960 -7420
rect 4800 -8260 5240 -7420
rect 6100 -8260 6540 -7420
rect 7380 -8260 7820 -7420
rect 8680 -8260 9120 -7420
rect 9940 -8260 10160 -7420
rect 3740 -8700 10180 -8260
rect 3740 -9540 3960 -8700
rect 4800 -9540 5240 -8700
rect 6100 -9540 6540 -8700
rect 7380 -9540 7820 -8700
rect 8680 -9540 9120 -8700
rect 9940 -9540 10160 -8700
rect 3740 -9840 10180 -9540
rect 3340 -17200 10180 -9840
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect 12600 -17200 13400 -16800
rect -9800 -17400 13400 -17200
rect -9800 -17800 -9200 -17400
rect 13000 -17800 13400 -17400
rect -9800 -18000 13400 -17800
<< viali >>
rect -9400 6200 13000 6600
rect -9600 -17000 -9200 5200
rect 4750 4995 5500 5045
rect -1488 4906 -1312 4940
rect -1168 4906 -992 4940
rect -1581 4710 -1547 4878
rect -933 4710 -899 4878
rect 1019 4710 1053 4878
rect -1488 4648 -1312 4682
rect -1168 4648 -992 4682
rect 1120 4400 1280 4440
rect -1500 4270 -1300 4304
rect -1140 4280 -1000 4340
rect -2300 4140 -2265 4205
rect -2242 4012 -1266 4046
rect 4360 4280 4400 4340
rect 4750 3995 5500 4045
rect -3200 3600 -2400 3800
rect 1120 3600 1280 3640
rect -1832 3260 -1772 3294
rect -1750 3055 -1715 3170
rect -1175 3025 -625 3075
rect -480 2860 -420 2960
rect 2160 2540 2220 2740
rect 5510 2690 5790 3460
rect 220 2220 260 2320
rect -480 1180 -420 1280
rect 220 800 260 1000
rect 2160 800 2220 1000
rect -1832 -16856 -1772 -16822
rect 2640 -2100 2780 -1620
rect 8560 -2080 8720 -1840
rect 1776 -7042 2890 -6645
rect 12800 -16800 13200 5400
rect -9200 -17800 13000 -17400
<< metal1 >>
rect -9800 6600 13400 6800
rect -9800 6200 -9400 6600
rect 13000 6200 13400 6600
rect -9800 6000 13400 6200
rect -9800 5200 -9000 6000
rect -9800 -17000 -9600 5200
rect -9200 -2080 -9000 5200
rect -2200 5120 6000 5640
rect 12600 5400 13400 6000
rect -2120 4560 -2040 5120
rect -1500 4940 -1300 5120
rect -1500 4906 -1488 4940
rect -1312 4906 -1300 4940
rect -1500 4900 -1300 4906
rect -1180 4940 -980 5120
rect -1180 4906 -1168 4940
rect -992 4906 -980 4940
rect -1180 4900 -980 4906
rect 1100 4900 1300 5120
rect 4740 5045 5530 5120
rect 4740 4995 4750 5045
rect 5500 4995 5530 5045
rect 4740 4980 5530 4995
rect -1587 4878 -1541 4890
rect -939 4880 -893 4890
rect -1587 4710 -1581 4878
rect -1547 4710 -1541 4878
rect -1587 4698 -1541 4710
rect -940 4878 1060 4880
rect -940 4710 -933 4878
rect -899 4710 1019 4878
rect 1053 4710 1060 4878
rect -940 4700 1060 4710
rect -939 4698 -893 4700
rect -1500 4682 -1300 4688
rect -1500 4630 -1490 4682
rect -1310 4630 -1300 4682
rect -1500 4620 -1300 4630
rect -1180 4682 -980 4688
rect -1180 4630 -1170 4682
rect -990 4630 -980 4682
rect -1180 4620 -980 4630
rect 1100 4630 1110 4680
rect 1290 4630 1300 4680
rect 1100 4620 1300 4630
rect -2120 4480 4240 4560
rect 1100 4442 1300 4450
rect 1100 4390 1120 4442
rect 1280 4390 1300 4442
rect -1180 4340 -980 4350
rect -1510 4330 -1290 4340
rect -1510 4320 -1500 4330
rect -1520 4270 -1500 4320
rect -1300 4320 -1290 4330
rect -1300 4270 -1280 4320
rect -1520 4260 -1280 4270
rect -1180 4280 -1140 4340
rect -1000 4280 -980 4340
rect -2325 4205 -2255 4220
rect -2325 4150 -2315 4205
rect -2260 4150 -2255 4205
rect -2325 4140 -2300 4150
rect -2265 4140 -2255 4150
rect -2325 4125 -2255 4140
rect -2255 4050 -1255 4055
rect -2260 4046 -1240 4050
rect -2260 4040 -2242 4046
rect -2620 4012 -2242 4040
rect -1266 4012 -1240 4046
rect -2620 3852 -1240 4012
rect -3332 3800 -1240 3852
rect -3332 3600 -3200 3800
rect -2400 3600 -1240 3800
rect -3332 3500 -1240 3600
rect -3332 3420 -2186 3500
rect -1180 3300 -980 4280
rect 1100 3640 1300 4390
rect 4160 3900 4240 4480
rect 4340 4340 4420 4360
rect 4400 4280 4420 4340
rect 4340 4260 4420 4280
rect 4720 4050 5520 4060
rect 4720 3995 4750 4050
rect 5500 3995 5520 4050
rect 4720 3980 5520 3995
rect 5840 3900 5920 5120
rect 4160 3820 5920 3900
rect 1100 3600 1120 3640
rect 1280 3600 1300 3640
rect 1100 3580 1300 3600
rect -1840 3294 -980 3300
rect -1840 3260 -1832 3294
rect -1772 3260 -980 3294
rect -1655 3185 -1610 3260
rect -1760 3170 -1610 3185
rect -1760 3055 -1750 3170
rect -1715 3155 -1610 3170
rect -1715 3055 -1705 3155
rect -1180 3140 -980 3260
rect 5480 3460 5860 3470
rect -1180 3100 -600 3140
rect -1760 3040 -1705 3055
rect -1200 3075 -600 3100
rect -1200 3025 -1175 3075
rect -625 3025 -600 3075
rect -1200 3000 -600 3025
rect -500 2960 -400 2980
rect -500 2860 -480 2960
rect -420 2860 -400 2960
rect -500 2840 -400 2860
rect 2140 2740 2240 2760
rect 2140 2540 2160 2740
rect 2220 2540 2240 2740
rect 5480 2690 5510 3460
rect 5790 2690 5860 3460
rect 5480 2650 5860 2690
rect 2140 2520 2240 2540
rect 200 2320 280 2340
rect 200 2220 220 2320
rect 200 2200 280 2220
rect -200 1700 500 1800
rect -200 1300 -60 1700
rect -500 1280 -60 1300
rect -500 1180 -480 1280
rect -420 1180 -60 1280
rect -500 1160 -60 1180
rect 200 1000 280 1020
rect 200 800 220 1000
rect 200 780 280 800
rect 2140 1000 2240 1020
rect 2140 800 2160 1000
rect 2220 800 2240 1000
rect 2140 780 2240 800
rect 480 -60 1960 140
rect -1440 -460 1960 -60
rect -9200 -17000 -2180 -2080
rect -9800 -17200 -2180 -17000
rect -1840 -16822 -1760 -16820
rect -1840 -16856 -1832 -16822
rect -1772 -16856 -1760 -16822
rect -1840 -17200 -1760 -16856
rect -1000 -17200 1200 -460
rect 2620 -1620 2800 -1600
rect 2620 -2100 2640 -1620
rect 2780 -2100 2800 -1620
rect 8540 -1840 8740 -1820
rect 8540 -2080 8560 -1840
rect 8720 -2080 8740 -1840
rect 8540 -2100 8740 -2080
rect 2620 -2120 2800 -2100
rect 4080 -4280 9860 -3660
rect 4080 -4960 4700 -4280
rect 5360 -4960 5980 -4280
rect 6660 -4960 7260 -4280
rect 7940 -4960 8560 -4280
rect 9240 -4960 9860 -4280
rect 4080 -5580 9860 -4960
rect 4080 -6630 4700 -5580
rect 1760 -6645 4700 -6630
rect 1760 -7042 1776 -6645
rect 2890 -7042 4700 -6645
rect 1760 -7060 4700 -7042
rect 4080 -7540 4700 -7060
rect 5360 -7540 5980 -5580
rect 7940 -7540 8560 -5580
rect 9240 -7540 9860 -5580
rect 4080 -8160 9860 -7540
rect 4080 -8820 4700 -8160
rect 5360 -8820 5980 -8160
rect 6660 -8820 7260 -8160
rect 7940 -8820 8560 -8160
rect 9240 -8820 9860 -8160
rect 4080 -9440 9860 -8820
rect 3740 -9840 10180 -9760
rect 3340 -17200 10180 -9840
rect 12600 -16800 12800 5400
rect 13200 -16800 13400 5400
rect 12600 -17200 13400 -16800
rect -9800 -17400 13400 -17200
rect -9800 -17800 -9200 -17400
rect 13000 -17800 13400 -17400
rect -9800 -18000 13400 -17800
<< via1 >>
rect -1490 4648 -1488 4682
rect -1488 4648 -1312 4682
rect -1312 4648 -1310 4682
rect -1490 4630 -1310 4648
rect -1170 4648 -1168 4682
rect -1168 4648 -992 4682
rect -992 4648 -990 4682
rect -1170 4630 -990 4648
rect 1110 4630 1290 4682
rect 1120 4440 1280 4442
rect 1120 4400 1280 4440
rect 1120 4390 1280 4400
rect -1500 4304 -1300 4330
rect -1500 4270 -1300 4304
rect -1140 4280 -1000 4340
rect -2315 4150 -2300 4205
rect -2300 4150 -2265 4205
rect -2265 4150 -2260 4205
rect 4340 4280 4360 4340
rect 4360 4280 4400 4340
rect 4750 4045 5500 4050
rect 4750 3995 5500 4045
rect -480 2860 -420 2960
rect 2160 2540 2220 2740
rect 5510 2690 5790 3460
rect 220 2220 260 2320
rect 260 2220 280 2320
rect 220 800 260 1000
rect 260 800 280 1000
rect 2160 800 2220 1000
rect 2640 -2100 2780 -1620
rect 8560 -2080 8720 -1840
rect 6740 -6700 7150 -6430
<< metal2 >>
rect -1500 4682 -1300 4690
rect -1500 4630 -1490 4682
rect -1310 4630 -1300 4682
rect -1500 4340 -1300 4630
rect -1180 4682 -980 4690
rect -1180 4630 -1170 4682
rect -990 4630 -980 4682
rect -1180 4360 -980 4630
rect 1100 4682 1300 4690
rect 1100 4630 1110 4682
rect 1290 4630 1300 4682
rect 1100 4442 1300 4630
rect 1100 4390 1120 4442
rect 1280 4390 1300 4442
rect -1180 4340 4400 4360
rect -1520 4330 -1280 4340
rect -1520 4270 -1500 4330
rect -1300 4270 -1280 4330
rect -1520 4260 -1280 4270
rect -1180 4280 -1140 4340
rect -1000 4280 4340 4340
rect -1180 4260 4400 4280
rect -2325 4205 -2255 4220
rect -2325 4150 -2315 4205
rect -2260 4200 -420 4205
rect -2260 4150 3680 4200
rect -2325 4140 3680 4150
rect -2325 4125 -2255 4140
rect -480 4080 3680 4140
rect -480 2980 -420 4080
rect 3540 3770 3680 4080
rect 4720 4050 5520 4060
rect 4720 3995 4750 4050
rect 5500 3995 5520 4050
rect 4720 3780 5520 3995
rect 4720 3770 5940 3780
rect 3540 3670 5940 3770
rect 5400 3460 5940 3670
rect -500 2960 -400 2980
rect -500 2860 -480 2960
rect -420 2860 -400 2960
rect -500 2840 -400 2860
rect 2140 2740 4380 2760
rect 2140 2540 2160 2740
rect 2220 2540 4380 2740
rect 2140 2520 4380 2540
rect 200 2320 2860 2340
rect 200 2220 220 2320
rect 280 2220 2860 2320
rect 200 2200 2860 2220
rect 180 1000 2240 1020
rect 180 800 220 1000
rect 280 800 2160 1000
rect 2220 800 2240 1000
rect 180 780 2240 800
rect 2540 -1620 2860 2200
rect 2540 -2100 2640 -1620
rect 2780 -2100 2860 -1620
rect 2540 -2240 2860 -2100
rect 3940 -1800 4380 2520
rect 5400 2690 5510 3460
rect 5790 2690 5940 3460
rect 5400 2460 5940 2690
rect 8500 -1800 9000 -1400
rect 3940 -1840 9000 -1800
rect 3940 -2080 8560 -1840
rect 8720 -2080 9000 -1840
rect 3940 -2140 9000 -2080
rect 8500 -6300 9000 -2140
rect 6700 -6430 9000 -6300
rect 6700 -6700 6740 -6430
rect 7150 -6700 9000 -6430
rect 6700 -6800 9000 -6700
use diff_pair  diff_pair_0
timestamp 1730311536
transform 1 0 -234 0 1 2300
box 234 -2300 2665 1550
use n20x1  n20x1_0
timestamp 1730304573
transform -1 0 -400 0 1 2600
box -100 -1200 1200 600
use n20x1  n20x1_1
timestamp 1730304573
transform -1 0 -400 0 1 1000
box -100 -1200 1200 600
use p20x05  p20x05_0
timestamp 1730605901
transform 1 0 1825 0 1 3470
box 2475 450 3975 1650
use sky130_fd_pr__nfet_01v8_6EEDFX  sky130_fd_pr__nfet_01v8_6EEDFX_0
timestamp 1730605901
transform 0 1 -1754 -1 0 4158
box -158 -526 158 526
use sky130_fd_pr__nfet_01v8_N7YW8T  sky130_fd_pr__nfet_01v8_N7YW8T_0
timestamp 1730605901
transform 0 1 -1802 -1 0 -1752
box -5058 -68 5058 68
use sky130_fd_pr__nfet_01v8_N7YW8T  sky130_fd_pr__nfet_01v8_N7YW8T_1
timestamp 1730605901
transform 0 1 -1802 -1 0 -11810
box -5058 -68 5058 68
use sky130_fd_pr__pfet_01v8_J24L55  sky130_fd_pr__pfet_01v8_J24L55_0
timestamp 1730316371
transform 0 1 1200 -1 0 4794
box -194 -200 194 200
use sky130_fd_pr__res_xhigh_po_5p73_G7V36E  sky130_fd_pr__res_xhigh_po_5p73_G7V36E_0
timestamp 1730605901
transform 1 0 2333 0 1 -4644
box -573 -2416 573 2416
use sky130_fd_pr__res_xhigh_po_5p73_QHLGXT  sky130_fd_pr__res_xhigh_po_5p73_QHLGXT_0
timestamp 1730605901
transform 1 0 -5243 0 1 2176
box -3057 -1676 3057 1676
use sky130_fd_pr__res_xhigh_po_5p73_QHLGXT  sky130_fd_pr__res_xhigh_po_5p73_QHLGXT_1
timestamp 1730605901
transform -1 0 -5243 0 1 -824
box -3057 -1676 3057 1676
use sky130_fd_pr__res_xhigh_po_5p73_QHLGXT  sky130_fd_pr__res_xhigh_po_5p73_QHLGXT_2
timestamp 1730605901
transform 0 1 7176 -1 0 557
box -3057 -1676 3057 1676
use sky130_fd_pr__res_xhigh_po_5p73_QHLGXT  sky130_fd_pr__res_xhigh_po_5p73_QHLGXT_3
timestamp 1730605901
transform 0 -1 4176 -1 0 557
box -3057 -1676 3057 1676
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 4 1288
timestamp 1730605901
transform 1 0 3716 0 1 -9796
box 0 0 1340 1340
<< labels >>
flabel metal1 200 5400 200 5400 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal2 5700 3700 5700 3700 0 FreeSans 1600 0 0 0 Vref
port 1 nsew
flabel viali -8200 -17600 -8200 -17600 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
<< end >>
