magic
tech sky130A
magscale 1 2
timestamp 1732923339
<< nwell >>
rect -194 -364 194 398
<< pmos >>
rect -100 -264 100 336
<< pdiff >>
rect -158 324 -100 336
rect -158 -252 -146 324
rect -112 -252 -100 324
rect -158 -264 -100 -252
rect 100 324 158 336
rect 100 -252 112 324
rect 146 -252 158 324
rect 100 -264 158 -252
<< pdiffc >>
rect -146 -252 -112 324
rect 112 -252 146 324
<< poly >>
rect -100 336 100 362
rect -100 -311 100 -264
rect -100 -345 -84 -311
rect 84 -345 100 -311
rect -100 -361 100 -345
<< polycont >>
rect -84 -345 84 -311
<< locali >>
rect -146 324 -112 340
rect -146 -268 -112 -252
rect 112 324 146 340
rect 112 -268 146 -252
rect -100 -345 -84 -311
rect 84 -345 100 -311
<< viali >>
rect -146 -252 -112 324
rect 112 -252 146 324
rect -84 -345 84 -311
<< metal1 >>
rect -152 324 -106 336
rect -152 -252 -146 324
rect -112 -252 -106 324
rect -152 -264 -106 -252
rect 106 324 152 336
rect 106 -252 112 324
rect 146 -252 152 324
rect 106 -264 152 -252
rect -96 -311 96 -305
rect -96 -345 -84 -311
rect 84 -345 96 -311
rect -96 -351 96 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__pfet_01v8_PXDZWB parameters
<< end >>
