magic
tech sky130A
magscale 1 2
timestamp 1731631080
<< xpolycontact >>
rect 131 1364 201 1796
rect -201 -1796 -131 -1364
<< xpolyres >>
rect -201 1190 35 1260
rect -201 -1364 -131 1190
rect -35 -1190 35 1190
rect 131 -1190 201 1364
rect -35 -1260 201 -1190
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 12.6 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 221.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string sky130_fd_pr__res_xhigh_po_0p35_BB2ZH9 parameters
<< end >>
